-- Entity name: modular_exponentiation_tb
-- Author: Luis Gallet, Jacob Barnett
-- Contact: luis.galletzambrano@mail.mcgill.ca, jacob.barnett@mail.mcgill.ca
-- Date: April 09, 2016
-- Description:

library ieee;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
--use IEEE.std_logic_arith.all;
--use IEEE.std_logic_unsigned.all;

entity modular_exponentiation_tb is
end entity;

architecture test of modular_exponentiation_tb is
-- define the ALU compontent to be tested
component modular_exponentiation is
 	generic(
		WIDTH_IN : integer := 512
	);
	port(	N :	in unsigned(WIDTH_IN-1 downto 0); --Number
		enc_dec : std_logic;
		--Exp :	in unsigned(WIDTH_IN-1 downto 0); --Exponent
		--M :	in unsigned(WIDTH_IN-1 downto 0); --Modulus
		--latch_in: in std_logic;
		clk :	in std_logic;
		reset :	in std_logic;
		C : 	out unsigned(WIDTH_IN-1 downto 0) --Output
		--C : out std_logic
	);

end component;

CONSTANT WIDTH_IN : integer := 512;

CONSTANT clk_period : time := 1 ns;

Signal M_in : unsigned(WIDTH_IN-1 downto 0) := (WIDTH_IN-1 downto 0 => '0');
Signal N_in : unsigned(WIDTH_IN-1 downto 0) := (WIDTH_IN-1 downto 0 => '0');
Signal Exp_in : unsigned(WIDTH_IN-1 downto 0) := (WIDTH_IN-1 downto 0 => '0');
signal latch_in : std_logic := '0';
signal enc_dec : std_logic;

Signal clk : std_logic := '0';
Signal reset_t : std_logic := '0';

Signal C_out : unsigned(WIDTH_IN-1 downto 0) := (WIDTH_IN-1 downto 0 => '0');
--signal c_out : std_logic;

Begin
-- device under test
dut: modular_exponentiation 
			generic map(WIDTH_IN => WIDTH_IN)
			PORT MAP(	N	=> 	N_in,
					enc_dec => 	enc_dec,
					--Exp 	=> 	Exp_in,
					--M 	=> 	M_in,
					--latch_in => latch_in,
					clk	=> 	clk,
					reset 	=>	reset_t,
					C	=>	C_out
				);
  
-- process for clock
clk_process : Process
Begin
	clk <= '0';
	wait for clk_period/2;
	clk <= '1';
	wait for clk_period/2;
end process;

stim_process: process
Begin


	reset_t <= '1';
	wait for 1 * clk_period;
	reset_t <= '0';
	wait for 1 * clk_period;


	REPORT "Begin test case for base=4446728192895187255737449916574481996753115952658605977007033762865282370651397068646324375752567034002689929313161372976205186035026701595623242884267844, exp=65537, mod=6874373683554289430325714128268458800697697146760798575501402831012475017846769541771555269176550565359325254833460767178884136299159177410149450184130651";
	REPORT "Expected output is 5126585062655550277416948279421250498005249302831876063220719451698168964783076608472238674806364148578582162270551448183956292595566138446551237116350418, 01100001111000100011100111001110011001001100110000100110010100101010111011111010100111001001011101010100011011100011001010000100100011011010110101011101010111100100000111110011100000101001111101101111011001101010100100100101100100110110111111011111010110111000110110011010001111010010010111101011000010000010000010111100000010010011101101110001101100111010010010000011010011101011100000101011001100010010000010100110001011110100110101011101100011001110001101010101100001101000000100111010111111001100111111010010";
	N_in <= "01010100111001110010011110010111000001001110010110011100001000001111110011010001101011110011001110001000111111110010100001010100001000111111110001110101111011001100000011011100100001100011000101101001011000100101110010100100110000101111110110111110111001100000001111011010100101110000011111011100001100010100000110101011110001000111110011010100010110101001111010100010110110101110011110100000000000011010100110010000010110100010100000101111010010011111100110010010101111010110101111010000001010010011111101000100";
	enc_dec <= '1';
	--Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	--M_in <= "10000011010000010011110100010110101100001100010010011111110101011001010111110100011000111101001110110100010101111110010110101001010000100101110110110011010111100111100001101010111001100011010001001001100001011011110101100000110011101001110010101101000100000011000100000111010000000001010000100101001011111111101010110100110011101100011000111011110100110001111010000101100000101010111110111001101100111110001001000111011101101110000111100100011010111000000011110110010110111000101111000111100100000000000001011011";
	wait for 526849 * clk_period;
	ASSERT(C_out = "01100001111000100011100111001110011001001100110000100110010100101010111011111010100111001001011101010100011011100011001010000100100011011010110101011101010111100100000111110011100000101001111101101111011001101010100100100101100100110110111111011111010110111000110110011010001111010010010111101011000010000010000010111100000010010011101101110001101100111010010010000011010011101011100000101011001100010010000010100110001011110100110101011101100011001110001101010101100001101000000100111010111111001100111111010010") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=5126585062655550277416948279421250498005249302831876063220719451698168964783076608472238674806364148578582162270551448183956292595566138446551237116350418, exp=1777412180414535825516414024192578762803034593464176447836661290133915026465475721791945195821650390919372264357709395823184803324327668922892527266987913, mod=6874373683554289430325714128268458800697697146760798575501402831012475017846769541771555269176550565359325254833460767178884136299159177410149450184130651";
	REPORT "Expected output is 4446728192895187255737449916574481996753115952658605977007033762865282370651397068646324375752567034002689929313161372976205186035026701595623242884267844, 01010100111001110010011110010111000001001110010110011100001000001111110011010001101011110011001110001000111111110010100001010100001000111111110001110101111011001100000011011100100001100011000101101001011000100101110010100100110000101111110110111110111001100000001111011010100101110000011111011100001100010100000110101011110001000111110011010100010110101001111010100010110110101110011110100000000000011010100110010000010110100010100000101111010010011111100110010010101111010110101111010000001010010011111101000100";
	N_in <= "01100001111000100011100111001110011001001100110000100110010100101010111011111010100111001001011101010100011011100011001010000100100011011010110101011101010111100100000111110011100000101001111101101111011001101010100100100101100100110110111111011111010110111000110110011010001111010010010111101011000010000010000010111100000010010011101101110001101100111010010010000011010011101011100000101011001100010010000010100110001011110100110101011101100011001110001101010101100001101000000100111010111111001100111111010010";
	enc_dec <= '0';
	--Exp_in <= "00100001111011111100111101001100101110111001110111001011001110011101110101010000110110000011001011010111110100010101011000110111010000100100101010011001111000110001011000111101100001011001001000000101011001001000100000000111101011001100010000010110100100011111010101111100011101111001100011001001101001100111111011101011010110110111011110011010011000100011100111100000111001001101001111011111100011101010000010011111010111101011101101010111001100100111000111011111101101011110010011001000111011000111111110001001";
	--M_in <= "10000011010000010011110100010110101100001100010010011111110101011001010111110100011000111101001110110100010101111110010110101001010000100101110110110011010111100111100001101010111001100011010001001001100001011011110101100000110011101001110010101101000100000011000100000111010000000001010000100101001011111111101010110100110011101100011000111011110100110001111010000101100000101010111110111001101100111110001001000111011101101110000111100100011010111000000011110110010110111000101111000111100100000000000001011011";
	wait for 526849 * clk_period;
	ASSERT(C_out = "01010100111001110010011110010111000001001110010110011100001000001111110011010001101011110011001110001000111111110010100001010100001000111111110001110101111011001100000011011100100001100011000101101001011000100101110010100100110000101111110110111110111001100000001111011010100101110000011111011100001100010100000110101011110001000111110011010100010110101001111010100010110110101110011110100000000000011010100110010000010110100010100000101111010010011111100110010010101111010110101111010000001010010011111101000100") REPORT "test failed" SEVERITY NOTE;




	wait;

end process;
end;

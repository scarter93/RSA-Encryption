-- Entity name: modular_exponentiation_tb
-- Author: Luis Gallet, Jacob Barnett
-- Contact: luis.galletzambrano@mail.mcgill.ca, jacob.barnett@mail.mcgill.ca
-- Date: April 07, 2016
-- Description:

library ieee;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
--use IEEE.std_logic_arith.all;
--use IEEE.std_logic_unsigned.all;

entity modular_exponentiation_tb is
end entity;

architecture test of modular_exponentiation_tb is
-- define the ALU compontent to be tested
component modular_exponentiation is
 	generic(
		WIDTH_IN : integer := 1024
	);
	port(	N :	in unsigned(WIDTH_IN-1 downto 0); --Number
		Exp :	in unsigned(WIDTH_IN-1 downto 0); --Exponent
		M :	in unsigned(WIDTH_IN-1 downto 0); --Modulus
		--latch_in: in std_logic;
		clk :	in std_logic;
		reset :	in std_logic;
		C : 	out unsigned(WIDTH_IN-1 downto 0) --Output
		--C : out std_logic
	);

end component;

CONSTANT WIDTH_IN : integer := 1024;

CONSTANT clk_period : time := 1 ns;

Signal M_in : unsigned(WIDTH_IN-1 downto 0) := (WIDTH_IN-1 downto 0 => '0');
Signal N_in : unsigned(WIDTH_IN-1 downto 0) := (WIDTH_IN-1 downto 0 => '0');
Signal Exp_in : unsigned(WIDTH_IN-1 downto 0) := (WIDTH_IN-1 downto 0 => '0');
signal latch_in : std_logic := '0';

Signal clk : std_logic := '0';
Signal reset_t : std_logic := '0';

Signal C_out : unsigned(WIDTH_IN-1 downto 0) := (WIDTH_IN-1 downto 0 => '0');
--signal c_out : std_logic;

Begin
-- device under test
dut: modular_exponentiation 
			generic map(WIDTH_IN => WIDTH_IN)
			PORT MAP(	N	=> 	N_in,
					Exp 	=> 	Exp_in,
					M 	=> 	M_in,
					--latch_in => latch_in,
					clk	=> 	clk,
					reset 	=>	reset_t,
					C	=>	C_out
				);
  
-- process for clock
clk_process : Process
Begin
	clk <= '0';
	wait for clk_period/2;
	clk <= '1';
	wait for clk_period/2;
end process;

stim_process: process
Begin


	reset_t <= '1';
	wait for 1 * clk_period;
	reset_t <= '0';
	wait for 1 * clk_period;

	REPORT "Begin test case for base=48710652365608707149836989914458686717733755910995547596578218050057100945316865280224526187143992460907135064440723548171898392370638635522044644519986320623387632295450866351690120114117289067800290142385269095764461988649384744426282338086430169792544780322814169332157155588941709143214823330323234993706, exp=65537, mod=101085849586972918373951121612216674320211056551798223901975548733952261029959998546313224140358869070834101471012517614081419683155460888808969783812042986057237910744195975198022337261915545878699256538888163262523218727463676472711933189488645397541286428123825701641111029164903115912968211727054649212211";
	REPORT "Expected output is 78799795239458298563353691390346558312549925708172243640699498939502899331534968131044595197610887613765223929325444718575462322694392030908519581712835019389768604995140350423198877676764850197073087744417715871071608677323963998156074041615272802459023814835942999844106835555664494494084023188374984383599, 0111000000110110111100100011010001001001101010001101111110110111110000001101000010011001100111110100011011000001010111001110010110011000011000101000000011111001100110110111111100110000111101000001101110101001001100000100101010011100100101010001010010110000010101001111010000010111111101001000000011111110011011000011100000011111111001001111000110101000011101011101111000001101101110000111010001000001110111101101110001010100010000110000001011000110101000000100011001110111011001011110010011100100100110111110101011001101000010000110110000110100111011110111001010000100101001011001011000011001000001101011011100111001011100000001001111100011010001110000000001101010000001101101110010111010000001110001001001010110111001100111101100100110110001111000010000001000110100010011000011100111110001100101110001010000110000110000100101111100011101100010111101110000100101000101111001000111101100111111010101110111110000110010111100101010100011100011100000111111100000000010111111010000111111000001011111111001011011001101110001101111";
	N_in <= "0100010101011101110000111111011111111000101010011000111010010011011100111101010111010001101011001001110110110010111100011100011111101000000011110000000001101110100110000000010011111110001101011110101111010101110011010001010011010000010011001010101011011011011010111111100101111111000111101101011110110111110110100111000100000101010011001111101010110001010010001010000000000011011111001011001110110001101110011101000000010101100101010111100011101110001100101111011001111100100011001101111101001011010001111100111101110001010011001011100101001011001011000011101110001011011010100111001010000010100100110101111111001011000001010011101000110110001101001100101011000010000000111111010100011000100110111011111011001100010100000010110000111010011000100000011000000111000000010100110100110100101100010110101000000010110110000101110111110000011001100100000001101111011100010100010101111110101001110000100010010011101100111101010011000010110010011010000111001101111111001010111000010110010111000010111100001111001100101011011000101010";
	Exp_in <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "1000111111110011011101101001001110010101100100101001001001101001111011001000100010110110101001000010001001110100011111110000100101101101111000100111111110101111001110011110001010000111001010011001001101101011011010111110111011011000101010100101011101001011100100000110010110010111110001110010011111110101001110110010001100100101010100011101001100001011100100101101001100111010010100101111101110010011000111101011000110000100010101100011001110000110100111001101110010101010110111101011111010100100100110100101111101101010110111111011101000110111100111111000110101011100011011110110101111111011101111000011101001010001011110000101011000100011101011001000110100100011110111010001111101000011110101000100101111011101001010110111110011000011001010100000000110001000110010111101000011001110010010001100010010101001111100001000001010100111101111001100101001010001010100010110100100000110000011001111110110011001110110010111110011101110101111101111100010010011010011101110010010100101101111110001010100100000110101001011110100110011";
	wait for 2102273 * clk_period;
	ASSERT(C_out = "0111000000110110111100100011010001001001101010001101111110110111110000001101000010011001100111110100011011000001010111001110010110011000011000101000000011111001100110110111111100110000111101000001101110101001001100000100101010011100100101010001010010110000010101001111010000010111111101001000000011111110011011000011100000011111111001001111000110101000011101011101111000001101101110000111010001000001110111101101110001010100010000110000001011000110101000000100011001110111011001011110010011100100100110111110101011001101000010000110110000110100111011110111001010000100101001011001011000011001000001101011011100111001011100000001001111100011010001110000000001101010000001101101110010111010000001110001001001010110111001100111101100100110110001111000010000001000110100010011000011100111110001100101110001010000110000110000100101111100011101100010111101110000100101000101111001000111101100111111010101110111110000110010111100101010100011100011100000111111100000000010111111010000111111000001011111111001011011001101110001101111") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=78799795239458298563353691390346558312549925708172243640699498939502899331534968131044595197610887613765223929325444718575462322694392030908519581712835019389768604995140350423198877676764850197073087744417715871071608677323963998156074041615272802459023814835942999844106835555664494494084023188374984383599, exp=56650153098712808734584689481872743861219031768839665646455558751554063248369178122419276076523193665160060405989711871614239011900663251662051066287667392590715022377626969748377874002370402201535558092016147265292815682771368956773202124425005250551323998958805203285195284823281515811871464589552798911681, mod=101085849586972918373951121612216674320211056551798223901975548733952261029959998546313224140358869070834101471012517614081419683155460888808969783812042986057237910744195975198022337261915545878699256538888163262523218727463676472711933189488645397541286428123825701641111029164903115912968211727054649212211";
	REPORT "Expected output is 48710652365608707149836989914458686717733755910995547596578218050057100945316865280224526187143992460907135064440723548171898392370638635522044644519986320623387632295450866351690120114117289067800290142385269095764461988649384744426282338086430169792544780322814169332157155588941709143214823330323234993706, 0100010101011101110000111111011111111000101010011000111010010011011100111101010111010001101011001001110110110010111100011100011111101000000011110000000001101110100110000000010011111110001101011110101111010101110011010001010011010000010011001010101011011011011010111111100101111111000111101101011110110111110110100111000100000101010011001111101010110001010010001010000000000011011111001011001110110001101110011101000000010101100101010111100011101110001100101111011001111100100011001101111101001011010001111100111101110001010011001011100101001011001011000011101110001011011010100111001010000010100100110101111111001011000001010011101000110110001101001100101011000010000000111111010100011000100110111011111011001100010100000010110000111010011000100000011000000111000000010100110100110100101100010110101000000010110110000101110111110000011001100100000001101111011100010100010101111110101001110000100010010011101100111101010011000010110010011010000111001101111111001010111000010110010111000010111100001111001100101011011000101010";
	N_in <= "0111000000110110111100100011010001001001101010001101111110110111110000001101000010011001100111110100011011000001010111001110010110011000011000101000000011111001100110110111111100110000111101000001101110101001001100000100101010011100100101010001010010110000010101001111010000010111111101001000000011111110011011000011100000011111111001001111000110101000011101011101111000001101101110000111010001000001110111101101110001010100010000110000001011000110101000000100011001110111011001011110010011100100100110111110101011001101000010000110110000110100111011110111001010000100101001011001011000011001000001101011011100111001011100000001001111100011010001110000000001101010000001101101110010111010000001110001001001010110111001100111101100100110110001111000010000001000110100010011000011100111110001100101110001010000110000110000100101111100011101100010111101110000100101000101111001000111101100111111010101110111110000110010111100101010100011100011100000111111100000000010111111010000111111000001011111111001011011001101110001101111";
	Exp_in <= "0101000010101100001010001010111111011101000010110001111101110010101011010101010010010000110001101011101101101000011111100010100101010010101000111011010011011011000001101001110110100101000100011110111111000100001010111110000011010111000110111101111110000000010000011001010000101101110100110011011011011001100000000010001011011010001011110101100100001111000010110110000111000101001101011110110000110111001011101110010001011101001111011101000111110010100001101100011001000100000110111101101111010010010000110101100101011001111000111010010100110001100111111010011010110100110001101000111110111011011010001101100100011110011101111011001101101001111011101111011100011010010111101111111001100101001111001001110010010000111110011111111110111010011110111111000100101100001001100100110010111101001010011001101001001000101100011001110000000001011011110000001000000111001010011101111111010010011010000111000101001101111010011011011101000001000001010100010111001111000101001011100110111000111011101001010010110010000010111100110011000001";
	M_in <= "1000111111110011011101101001001110010101100100101001001001101001111011001000100010110110101001000010001001110100011111110000100101101101111000100111111110101111001110011110001010000111001010011001001101101011011010111110111011011000101010100101011101001011100100000110010110010111110001110010011111110101001110110010001100100101010100011101001100001011100100101101001100111010010100101111101110010011000111101011000110000100010101100011001110000110100111001101110010101010110111101011111010100100100110100101111101101010110111111011101000110111100111111000110101011100011011110110101111111011101111000011101001010001011110000101011000100011101011001000110100100011110111010001111101000011110101000100101111011101001010110111110011000011001010100000000110001000110010111101000011001110010010001100010010101001111100001000001010100111101111001100101001010001010100010110100100000110000011001111110110011001110110010111110011101110101111101111100010010011010011101110010010100101101111110001010100100000110101001011110100110011";
	wait for 2102273 * clk_period;
	ASSERT(C_out = "0100010101011101110000111111011111111000101010011000111010010011011100111101010111010001101011001001110110110010111100011100011111101000000011110000000001101110100110000000010011111110001101011110101111010101110011010001010011010000010011001010101011011011011010111111100101111111000111101101011110110111110110100111000100000101010011001111101010110001010010001010000000000011011111001011001110110001101110011101000000010101100101010111100011101110001100101111011001111100100011001101111101001011010001111100111101110001010011001011100101001011001011000011101110001011011010100111001010000010100100110101111111001011000001010011101000110110001101001100101011000010000000111111010100011000100110111011111011001100010100000010110000111010011000100000011000000111000000010100110100110100101100010110101000000010110110000101110111110000011001100100000001101111011100010100010101111110101001110000100010010011101100111101010011000010110010011010000111001101111111001010111000010110010111000010111100001111001100101011011000101010") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=52945756746696132404706099581856910543193155207381989436042422850102363321984001351876898590441763010659051864378460269214251602217399703843165383350575434618971818324841503807764858686740007010189230709233762922734409247777204723056980424707153048058553912823586297528936634788155150929443130274883441810018, exp=65537, mod=91614999902063619993535257798090717108166556845768742750053702671887332260227750111395462504643993758854755991446422864968374522909645384275889871099632510981745375395280657289104997539222681158988688440764880230613021164250551518766136363464492794503234577373221231297820270229024966220822597694881823728601";
	REPORT "Expected output is 50015781274980223515381148350956242357843833061531049273321924445588310457485306214614429816636744925046308628508957997208771448718659888849560772086041276716811447444300656099521114306850442419482313227481118639104445234349627131260592028106646784400849249488688111098761385743107871265071715488296427609782, 0100011100111001100011101110011011001000011001100101100011010001110000110101111111110100110010011011111111110001001100110001101110011000010001111001001110010111010110110011101011001111110000000001110110010100001100011100111110011011111110100001101110000011010100101100100011111010100011111000110010101111010100101111011000010100111000100100101000010101101100111011000111011100110000110001110110110011010001100100010100011110011001010111001011001001010011100000000111100101100110010110100001110111101110101000011000010000100110000111111011101110110000111111111100101101111100001101001111101100101111000111110110011011001110010011010001010010001011110011111100110001111110000011001110100000001101001110101100011010111010010100001011100000010010111010010111011011100101111010101111010010000000001011101011000011010011000111011110010100111100110000010001110111101010011001100001000011001011110111100011100011111100110010000110010001011100000100011000011000000011111101001111011101100011001110010011110100111000000101111010110110";
	N_in <= "0100101101100101101100101101101001000010110001000101111010111001011001010100001001100011111011100100001110101110001110110011011001000101001010010000011111110010111010000000001110010000101100111011011100111010101110010101011110111001000100110010111010010110001010011100001110010001001011110001101010100111111101101001110000101101111000000000011100010010100101110111100101011110111001111100000000010001001011010011000010110000011111011010111101101010100010010010001110101000101110000001001111100100101011111000110111000100101010101101001110100100101110100111011101101001011010110001110110000100001011000001101000110011111000000100111011011001011101010010111101100110111001100110000110101100100011001001001100000101101000000110011110000100110001000001100111011101011101111110111000010000111010110001011111100100010110000111001100111100011001011000010101110110100000011110101100010011100111000110000000110111101100011001101111111110010111001101001110100111011100101110101011111110110110101010111001010001011000000101101001100010";
	Exp_in <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "1000001001110110110011101010000110111100001001100111000101100100000000101101011001000101101010000100001101111111101011001010100110110110000010101111101011001100011010000101001000111010110101110000111011001101100011000111001000110110101111101000001000000001001101101001101100101100000100101010011111001011111110101100101101111011000110100001110110110000001100010010110110011010110011110000110100101011110101010100100100010011111010101000010101000111100111010101011010111100011000010101111111111111110111001100001100001011111111100111100011100110101010000001000010001010100101110101001111111010100001011011111011100100001101011001100111111000011111000001110100110011101100001010110000110100010010110110001000110001111000101001000010011111000010110111001011100100110011010100000011101000010111000101100010100001111101101010010100111111000101001111010000001110100111111110001100000110110100000101101110010110000001110111101011010101011000111101000110010101011011001000110011111100010001100111010101011101110001000010001111011001";
	wait for 2102273 * clk_period;
	ASSERT(C_out = "0100011100111001100011101110011011001000011001100101100011010001110000110101111111110100110010011011111111110001001100110001101110011000010001111001001110010111010110110011101011001111110000000001110110010100001100011100111110011011111110100001101110000011010100101100100011111010100011111000110010101111010100101111011000010100111000100100101000010101101100111011000111011100110000110001110110110011010001100100010100011110011001010111001011001001010011100000000111100101100110010110100001110111101110101000011000010000100110000111111011101110110000111111111100101101111100001101001111101100101111000111110110011011001110010011010001010010001011110011111100110001111110000011001110100000001101001110101100011010111010010100001011100000010010111010010111011011100101111010101111010010000000001011101011000011010011000111011110010100111100110000010001110111101010011001100001000011001011110111100011100011111100110010000110010001011100000100011000011000000011111101001111011101100011001110010011110100111000000101111010110110") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=50015781274980223515381148350956242357843833061531049273321924445588310457485306214614429816636744925046308628508957997208771448718659888849560772086041276716811447444300656099521114306850442419482313227481118639104445234349627131260592028106646784400849249488688111098761385743107871265071715488296427609782, exp=6742132604904906224404848381222691435565975001405963749996322809809918114821832534099215949156933974685391277396678173821543102735755675242422091942859931797281878310870139536224340338415724312865283362257014161613435849987783434968713772954266748032566615144404623338638208093287338958227687842861645180973, mod=91614999902063619993535257798090717108166556845768742750053702671887332260227750111395462504643993758854755991446422864968374522909645384275889871099632510981745375395280657289104997539222681158988688440764880230613021164250551518766136363464492794503234577373221231297820270229024966220822597694881823728601";
	REPORT "Expected output is 52945756746696132404706099581856910543193155207381989436042422850102363321984001351876898590441763010659051864378460269214251602217399703843165383350575434618971818324841503807764858686740007010189230709233762922734409247777204723056980424707153048058553912823586297528936634788155150929443130274883441810018, 0100101101100101101100101101101001000010110001000101111010111001011001010100001001100011111011100100001110101110001110110011011001000101001010010000011111110010111010000000001110010000101100111011011100111010101110010101011110111001000100110010111010010110001010011100001110010001001011110001101010100111111101101001110000101101111000000000011100010010100101110111100101011110111001111100000000010001001011010011000010110000011111011010111101101010100010010010001110101000101110000001001111100100101011111000110111000100101010101101001110100100101110100111011101101001011010110001110110000100001011000001101000110011111000000100111011011001011101010010111101100110111001100110000110101100100011001001001100000101101000000110011110000100110001000001100111011101011101111110111000010000111010110001011111100100010110000111001100111100011001011000010101110110100000011110101100010011100111000110000000110111101100011001101111111110010111001101001110100111011100101110101011111110110110101010111001010001011000000101101001100010";
	N_in <= "0100011100111001100011101110011011001000011001100101100011010001110000110101111111110100110010011011111111110001001100110001101110011000010001111001001110010111010110110011101011001111110000000001110110010100001100011100111110011011111110100001101110000011010100101100100011111010100011111000110010101111010100101111011000010100111000100100101000010101101100111011000111011100110000110001110110110011010001100100010100011110011001010111001011001001010011100000000111100101100110010110100001110111101110101000011000010000100110000111111011101110110000111111111100101101111100001101001111101100101111000111110110011011001110010011010001010010001011110011111100110001111110000011001110100000001101001110101100011010111010010100001011100000010010111010010111011011100101111010101111010010000000001011101011000011010011000111011110010100111100110000010001110111101010011001100001000011001011110111100011100011111100110010000110010001011100000100011000011000000011111101001111011101100011001110010011110100111000000101111010110110";
	Exp_in <= "0000100110011001111000101011010100000110010110101011000111100111100100010100100111100001100100000111001101111111001101101101111010111010011101011110111001100101000100101001110001010010100101100011011100010001101010110110111101010000010101100000111011001101001101100000111010001111010111001100010000011010011111111101011101101111101101001100100101010000100010010001110111111001000100011001100110111111100010110000111110111000101101100111111010011110011110011001011011000011100000000011110011100000000010000001111000010010010110111111100111011101101001100010100110011110101100000000100101010001101111011010011110010100100110101101011000101000100110001011011001100111100101110001011110011111111111001010101011111011101110100010010111001011101101101101111011100110111000010101010100111100011111100110111110000111010110111000100101011111000011111111101001100000100011011111101001111100010010110010000010111010111100111001001101110101001011101101011011100010111100011110001001110101101110000101010010101000000100100011000000101101";
	M_in <= "1000001001110110110011101010000110111100001001100111000101100100000000101101011001000101101010000100001101111111101011001010100110110110000010101111101011001100011010000101001000111010110101110000111011001101100011000111001000110110101111101000001000000001001101101001101100101100000100101010011111001011111110101100101101111011000110100001110110110000001100010010110110011010110011110000110100101011110101010100100100010011111010101000010101000111100111010101011010111100011000010101111111111111110111001100001100001011111111100111100011100110101010000001000010001010100101110101001111111010100001011011111011100100001101011001100111111000011111000001110100110011101100001010110000110100010010110110001000110001111000101001000010011111000010110111001011100100110011010100000011101000010111000101100010100001111101101010010100111111000101001111010000001110100111111110001100000110110100000101101110010110000001110111101011010101011000111101000110010101011011001000110011111100010001100111010101011101110001000010001111011001";
	wait for 2102273 * clk_period;
	ASSERT(C_out = "0100101101100101101100101101101001000010110001000101111010111001011001010100001001100011111011100100001110101110001110110011011001000101001010010000011111110010111010000000001110010000101100111011011100111010101110010101011110111001000100110010111010010110001010011100001110010001001011110001101010100111111101101001110000101101111000000000011100010010100101110111100101011110111001111100000000010001001011010011000010110000011111011010111101101010100010010010001110101000101110000001001111100100101011111000110111000100101010101101001110100100101110100111011101101001011010110001110110000100001011000001101000110011111000000100111011011001011101010010111101100110111001100110000110101100100011001001001100000101101000000110011110000100110001000001100111011101011101111110111000010000111010110001011111100100010110000111001100111100011001011000010101110110100000011110101100010011100111000110000000110111101100011001101111111110010111001101001110100111011100101110101011111110110110101010111001010001011000000101101001100010") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=63458902791780287686094709450925892091127662722534075683020607787091115978366520003136195452962212645585642620691088135044662624633457008091771095535465805863596317316685108194400452046939069656769732272945471594014223928009546113760330098159915441574673773583938261815164965977033033424030068706240845418333, exp=65537, mod=93913334683773701655465005322140809550548642280383822567732640479866935892980619197652902575692747797499373133459790026848425700563099723476455918470997530928429009082187450219255838985189723601331723477898566474599953344750767563740779093354894961458592293472647658095410540308249818616262852063442988090421";
	REPORT "Expected output is 21895668108373993532791060793102974360094722833748931149563219520266259367088222909192512775549108764775036770718118410699487113818360708481886898244139698963085114998360260980824720905707677678859241758663616182106970266406425915700221725335727049860217679918083837457415561437852386831984812405273303966650, 0001111100101110001100110000101101111010011010100110011011000101010101101100100011001010010110000010001000101001001110000000011111000011100111100101101000101110111111100101001000111110111100100110001110010111001000110011100000110010111001011111000000100001100011110100010111001100100001010000111010010000111010000101100011101111111001101111100110000101010001100101000111111111101110100100100110101000000001100101000100100111111010100000100101011110110100010100101010001111111011010110111110000011001000011001000110100100101101011111000001101000010100001100100011011111111111100101010111100001010000000000001101100101011101111010001101100010001010011100000001101001011111111101001011111101111101101101100100001000110011110011000100111000101011001010111110111001111010101111011011011001100010100110110111010010010100100010101001111010101110000111000110010110011100011001100101101111101000001011100110110111011111000001101001011111100110001110101010011001101100010100011010001010100110100101110111100100101011111110001110111010";
	N_in <= "0101101001011110010101001000011001001010001110011011000010101000111001011111101000101111100001000111010100110011111010100111111010000010010010111010100001100000010110101101100011010111110111101100101110111001000100100010100000111111011100010000111001011100001101101000111010001111000001001011100100110010011011111111011011110101111000001010111000010100110111010111010010001110011010101011000001101000100010101100111111001010000011000010111100000111000100110111100000100011110101100010011101011111010101101001101001000000011111000001001001111001111110111101011000010000010011101101011010110101011111110111010111101011010010110011101010000110001101100001011110111111001011110111111001000001111001000000001010111110111010000101011100101000001101000111011100001011000000100100011100011101101001100010100111110000001010011001101001110000110110000000100101000001000100111010111010010011110011111100011111011000000010110110101111111010101000101100101100101001011110001000111011011001011001101010100010000111001010011000111101011101";
	Exp_in <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "1000010110111100101011011101101011110010110111000010100001011010001010010010111000010000111001110110101101001011011000011011000010101010010010011100110111100111011100111101110001101011000110110100010010000010100101111100000110000000000111111011001010101010011110110010011011000000001001000001101010011011111111010011001000110011011111010000111100011011001011110001010100111101010011101000101011000011001001010001100111101011110001010101111101101001011010100101000000000001100000101111100000011010110100011101001111011010011000111010001001010010101100001100011100010001111100111100011010000100001000100111101000001011010100011010011100000101111110100101010110001110000011000010100111110110111111011100000010110101001110110010000001111011110010010000111001010010111100010111011111111101111110001110011101111110101110111110000001101001101000001001010101111101011000001010101100010000011001110010010101001000100111001111011101001010100010001000011110100100011010111010100011100000010101011100001111111000101111101100010000110101";
	wait for 2102273 * clk_period;
	ASSERT(C_out = "0001111100101110001100110000101101111010011010100110011011000101010101101100100011001010010110000010001000101001001110000000011111000011100111100101101000101110111111100101001000111110111100100110001110010111001000110011100000110010111001011111000000100001100011110100010111001100100001010000111010010000111010000101100011101111111001101111100110000101010001100101000111111111101110100100100110101000000001100101000100100111111010100000100101011110110100010100101010001111111011010110111110000011001000011001000110100100101101011111000001101000010100001100100011011111111111100101010111100001010000000000001101100101011101111010001101100010001010011100000001101001011111111101001011111101111101101101100100001000110011110011000100111000101011001010111110111001111010101111011011011001100010100110110111010010010100100010101001111010101110000111000110010110011100011001100101101111101000001011100110110111011111000001101001011111100110001110101010011001101100010100011010001010100110100101110111100100101011111110001110111010") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=21895668108373993532791060793102974360094722833748931149563219520266259367088222909192512775549108764775036770718118410699487113818360708481886898244139698963085114998360260980824720905707677678859241758663616182106970266406425915700221725335727049860217679918083837457415561437852386831984812405273303966650, exp=83719101457651570438336085050207249589875998717470498586670797484707356083977092564268665443637905375182047951174471103934656372797015047143826871357321434267260677763431640642220794773402049979704338225738604453723814317468090945660854650170656389489765272399565922785628859204050572994478716811050334621473, mod=93913334683773701655465005322140809550548642280383822567732640479866935892980619197652902575692747797499373133459790026848425700563099723476455918470997530928429009082187450219255838985189723601331723477898566474599953344750767563740779093354894961458592293472647658095410540308249818616262852063442988090421";
	REPORT "Expected output is 63458902791780287686094709450925892091127662722534075683020607787091115978366520003136195452962212645585642620691088135044662624633457008091771095535465805863596317316685108194400452046939069656769732272945471594014223928009546113760330098159915441574673773583938261815164965977033033424030068706240845418333, 0101101001011110010101001000011001001010001110011011000010101000111001011111101000101111100001000111010100110011111010100111111010000010010010111010100001100000010110101101100011010111110111101100101110111001000100100010100000111111011100010000111001011100001101101000111010001111000001001011100100110010011011111111011011110101111000001010111000010100110111010111010010001110011010101011000001101000100010101100111111001010000011000010111100000111000100110111100000100011110101100010011101011111010101101001101001000000011111000001001001111001111110111101011000010000010011101101011010110101011111110111010111101011010010110011101010000110001101100001011110111111001011110111111001000001111001000000001010111110111010000101011100101000001101000111011100001011000000100100011100011101101001100010100111110000001010011001101001110000110110000000100101000001000100111010111010010011110011111100011111011000000010110110101111111010101000101100101100101001011110001000111011011001011001101010100010000111001010011000111101011101";
	N_in <= "0001111100101110001100110000101101111010011010100110011011000101010101101100100011001010010110000010001000101001001110000000011111000011100111100101101000101110111111100101001000111110111100100110001110010111001000110011100000110010111001011111000000100001100011110100010111001100100001010000111010010000111010000101100011101111111001101111100110000101010001100101000111111111101110100100100110101000000001100101000100100111111010100000100101011110110100010100101010001111111011010110111110000011001000011001000110100100101101011111000001101000010100001100100011011111111111100101010111100001010000000000001101100101011101111010001101100010001010011100000001101001011111111101001011111101111101101101100100001000110011110011000100111000101011001010111110111001111010101111011011011001100010100110110111010010010100100010101001111010101110000111000110010110011100011001100101101111101000001011100110110111011111000001101001011111100110001110101010011001101100010100011010001010100110100101110111100100101011111110001110111010";
	Exp_in <= "0111011100111000010011110010100000001011001011100011011000001110110000011111110100011101111101101001111101010000100100001110001011000011101110111000110110000001110100100110100001100001010101101110101010001001000111001010110111010100000000001110110111101110010010100110000010101110000100101100000101100001111000111010001000111000000000100011100101010000001110110111010111001100101101000101001011000001010010100011011011000100010101101010110000001010101101100100101001100010001111011110111100111000001001110110110000100000010000110111000101101000001010011011110101101100100001001001001101110010000110000110100111100000101111010010100000110111111010101011110100001011101101101101011111011010110010001000110010111110010111000100001011100110111101111001011011111111100111000001011000000001010111001011101110001100001111101101111000010101010011110010001000000010111010000011000000010100101001000100001111110000000101111011000110000101000111000110010111100011101011010001100011011011001101110110100100111100001111010000111100100001";
	M_in <= "1000010110111100101011011101101011110010110111000010100001011010001010010010111000010000111001110110101101001011011000011011000010101010010010011100110111100111011100111101110001101011000110110100010010000010100101111100000110000000000111111011001010101010011110110010011011000000001001000001101010011011111111010011001000110011011111010000111100011011001011110001010100111101010011101000101011000011001001010001100111101011110001010101111101101001011010100101000000000001100000101111100000011010110100011101001111011010011000111010001001010010101100001100011100010001111100111100011010000100001000100111101000001011010100011010011100000101111110100101010110001110000011000010100111110110111111011100000010110101001110110010000001111011110010010000111001010010111100010111011111111101111110001110011101111110101110111110000001101001101000001001010101111101011000001010101100010000011001110010010101001000100111001111011101001010100010001000011110100100011010111010100011100000010101011100001111111000101111101100010000110101";
	wait for 2102273 * clk_period;
	ASSERT(C_out = "0101101001011110010101001000011001001010001110011011000010101000111001011111101000101111100001000111010100110011111010100111111010000010010010111010100001100000010110101101100011010111110111101100101110111001000100100010100000111111011100010000111001011100001101101000111010001111000001001011100100110010011011111111011011110101111000001010111000010100110111010111010010001110011010101011000001101000100010101100111111001010000011000010111100000111000100110111100000100011110101100010011101011111010101101001101001000000011111000001001001111001111110111101011000010000010011101101011010110101011111110111010111101011010010110011101010000110001101100001011110111111001011110111111001000001111001000000001010111110111010000101011100101000001101000111011100001011000000100100011100011101101001100010100111110000001010011001101001110000110110000000100101000001000100111010111010010011110011111100011111011000000010110110101111111010101000101100101100101001011110001000111011011001011001101010100010000111001010011000111101011101") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=86839933975437002323963202225608757216981170417209756336946833671590005618973644873486967270266117361008160186582025163334060833773022340084139943422622102813746160832541702585141883794218254222340773583261983690741376470958298461709208863065882912105823635366194326115616517079719314203121092710944896792856, exp=65537, mod=146367340704051091293657330190128348760950155057778814316980525199527483741156987495468650741297321347767126517041298280090821875685866758748325900594251354037522736860962097760695802601558720999885522619682101995810565712896793382735322184664507538870977581576818286890910286020450716192664810991677323322149";
	REPORT "Expected output is 132533347433158961750583937752889294979220196163280066140789635676495940178544157436631797453762693836241835968670015021814572444650187204063490617063281058672642120548448685886013691815936055492528466462305411906079059876385312790244119941527897272274104375119172750702797656694883181920222855503365527744074, 1011110010111011110101110010001111001000101101110001111110101000101011101001010001000010111000110001111011110110110110101100101111000101010111101110001000010000010011111010011101000111010010011111101001011001110111110010001110001000101011110000001101000010011100101001101101001010101010010101100111111100101001101001110001001011010101001111100111000110100100101100000011010101000011111111010100000100011000100111110100111010101010010111110111111011001001101110010110001101010001101001100111010111110100100111100011101101110110100001101100010111111111100001001000000110010000011001110101000101110110000111101001101101000101100010110100111101010010111010001000000000000000011101001011011110000101101101011100000101111011100101111000000000100111001100010011001000000001101001000101110010010000110010101110000010010100010100101000101010110001010001011011101101100010101001000010000110010100010111111101111110101011101010111110101011110110100111111011100010100101100110000101011011101000110011101100000011001001101010111001001010";
	N_in <= "0111101110101010000001110001100111101011100000000000001010001001001100110100000110011110001000110000001000100000011100100101110010010110110010110011000000011100001100010011110100111001000011010001010101101010111110011011111100000110010101111000011010101001000101011101011111011111110011001011010101000011010001010110000110011001010110101010000100110111001100001110101111000011111111111011000011101000011011101100000101010100100111101011011101110101111010010011010101001001101000010000111111010001111111001000001100111011110010000101001111111010101011000110110110000101001101000111000000011111000110010000110111101000101011111110101111001001001000100010110100010110000011110000100010000101010110111111000011001101001100011111110010111011110000110000000011000000110011110000010000001000101110000110010000000110100111110110001100010001111111011001001010000011110011101000001011000101010111000000111110001010010101000101110101110101110000011011010001101111000010101011010110010110100001011111000101110010100000010011100100011000";
	Exp_in <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "1101000001101111000110110110011011010000010010000000000010000111100101101111101100000011100110011100110011011011110100010110001010010101111111100001101111010110011111000001000001011000100000101011101000111100010110110101000101100011000001001010110111010101111100001100110100011110110000011100101000100100010101001111000111111101111011010110010111100001011111001010010001011110101001110111010100111100101001110110001101000100101010010100001001000110111011000000100110110101001001011000100101101010011110010010000000110100000110110011011110111111011100111100001100001000101011111010011001111000010100000011100101001011111000000001110000111101101010100100010100001010101110001011000100101010110100000110011000110101001010001000010110001010010110000100011100010111101000101001010111000010110101011100111100101110101110010111010111110101011001000011011101001101110111010100011011110111000100001000001100001110010111011011010100010010110000100000101000110100100111000110100010100000011010100000101001111010000001111010001100100101";
	wait for 2102273 * clk_period;
	ASSERT(C_out = "1011110010111011110101110010001111001000101101110001111110101000101011101001010001000010111000110001111011110110110110101100101111000101010111101110001000010000010011111010011101000111010010011111101001011001110111110010001110001000101011110000001101000010011100101001101101001010101010010101100111111100101001101001110001001011010101001111100111000110100100101100000011010101000011111111010100000100011000100111110100111010101010010111110111111011001001101110010110001101010001101001100111010111110100100111100011101101110110100001101100010111111111100001001000000110010000011001110101000101110110000111101001101101000101100010110100111101010010111010001000000000000000011101001011011110000101101101011100000101111011100101111000000000100111001100010011001000000001101001000101110010010000110010101110000010010100010100101000101010110001010001011011101101100010101001000010000110010100010111111101111110101011101010111110101011110110100111111011100010100101100110000101011011101000110011101100000011001001101010111001001010") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=132533347433158961750583937752889294979220196163280066140789635676495940178544157436631797453762693836241835968670015021814572444650187204063490617063281058672642120548448685886013691815936055492528466462305411906079059876385312790244119941527897272274104375119172750702797656694883181920222855503365527744074, exp=79489546215703899191660461969987155181038770752650618111448050000787069919515075437366986849935979086771252376436728693486008395248659073155170566596417812668987475554333258389924103505907986063479536767056114802597237522843783921675869122149426399735079325720999564892573278117471627648045327170749357047393, mod=146367340704051091293657330190128348760950155057778814316980525199527483741156987495468650741297321347767126517041298280090821875685866758748325900594251354037522736860962097760695802601558720999885522619682101995810565712896793382735322184664507538870977581576818286890910286020450716192664810991677323322149";
	REPORT "Expected output is 86839933975437002323963202225608757216981170417209756336946833671590005618973644873486967270266117361008160186582025163334060833773022340084139943422622102813746160832541702585141883794218254222340773583261983690741376470958298461709208863065882912105823635366194326115616517079719314203121092710944896792856, 0111101110101010000001110001100111101011100000000000001010001001001100110100000110011110001000110000001000100000011100100101110010010110110010110011000000011100001100010011110100111001000011010001010101101010111110011011111100000110010101111000011010101001000101011101011111011111110011001011010101000011010001010110000110011001010110101010000100110111001100001110101111000011111111111011000011101000011011101100000101010100100111101011011101110101111010010011010101001001101000010000111111010001111111001000001100111011110010000101001111111010101011000110110110000101001101000111000000011111000110010000110111101000101011111110101111001001001000100010110100010110000011110000100010000101010110111111000011001101001100011111110010111011110000110000000011000000110011110000010000001000101110000110010000000110100111110110001100010001111111011001001010000011110011101000001011000101010111000000111110001010010101000101110101110101110000011011010001101111000010101011010110010110100001011111000101110010100000010011100100011000";
	N_in <= "1011110010111011110101110010001111001000101101110001111110101000101011101001010001000010111000110001111011110110110110101100101111000101010111101110001000010000010011111010011101000111010010011111101001011001110111110010001110001000101011110000001101000010011100101001101101001010101010010101100111111100101001101001110001001011010101001111100111000110100100101100000011010101000011111111010100000100011000100111110100111010101010010111110111111011001001101110010110001101010001101001100111010111110100100111100011101101110110100001101100010111111111100001001000000110010000011001110101000101110110000111101001101101000101100010110100111101010010111010001000000000000000011101001011011110000101101101011100000101111011100101111000000000100111001100010011001000000001101001000101110010010000110010101110000010010100010100101000101010110001010001011011101101100010101001000010000110010100010111111101111110101011101010111110101011110110100111111011100010100101100110000101011011101000110011101100000011001001101010111001001010";
	Exp_in <= "0111000100110010011001100010011101001000001001100101001001100011010100001101001110110001111110001110110100010000110101000111111000111110000001110110101100000110111010010000100111010111100001111110011110101100101011111100101101011011100000110100011100000101010100010110100110010100101100101001101000011101011100010010010010011011010010110011101001110001011000110100011111000001010000000010000010100011011110000010010010101001001111010110001100001001001100010101011101110100010100010000110010110100011111101101010101111011110011111010101101101110100101000011100001111100110000101001000000111000000101101111100100110110111000000111110110111101001110111001110100010100011001101110001111010001011110001111100011001000011010000111000010110100001110110011011000000111000111100101001011111101110001110010100101001100100010001111101100000001010000111001100011010110001011000000110001110101101101001110100000100111011101000111001100101001010001010001011010011100010101101111100010101100111000100100101110000100111001110011111001100001";
	M_in <= "1101000001101111000110110110011011010000010010000000000010000111100101101111101100000011100110011100110011011011110100010110001010010101111111100001101111010110011111000001000001011000100000101011101000111100010110110101000101100011000001001010110111010101111100001100110100011110110000011100101000100100010101001111000111111101111011010110010111100001011111001010010001011110101001110111010100111100101001110110001101000100101010010100001001000110111011000000100110110101001001011000100101101010011110010010000000110100000110110011011110111111011100111100001100001000101011111010011001111000010100000011100101001011111000000001110000111101101010100100010100001010101110001011000100101010110100000110011000110101001010001000010110001010010110000100011100010111101000101001010111000010110101011100111100101110101110010111010111110101011001000011011101001101110111010100011011110111000100001000001100001110010111011011010100010010110000100000101000110100100111000110100010100000011010100000101001111010000001111010001100100101";
	wait for 2102273 * clk_period;
	ASSERT(C_out = "0111101110101010000001110001100111101011100000000000001010001001001100110100000110011110001000110000001000100000011100100101110010010110110010110011000000011100001100010011110100111001000011010001010101101010111110011011111100000110010101111000011010101001000101011101011111011111110011001011010101000011010001010110000110011001010110101010000100110111001100001110101111000011111111111011000011101000011011101100000101010100100111101011011101110101111010010011010101001001101000010000111111010001111111001000001100111011110010000101001111111010101011000110110110000101001101000111000000011111000110010000110111101000101011111110101111001001001000100010110100010110000011110000100010000101010110111111000011001101001100011111110010111011110000110000000011000000110011110000010000001000101110000110010000000110100111110110001100010001111111011001001010000011110011101000001011000101010111000000111110001010010101000101110101110101110000011011010001101111000010101011010110010110100001011111000101110010100000010011100100011000") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=54051473182883694870366764758765700911582559777313054613910121608584026737001907012426262195401178256691273833725480698483655594641432143815158493354852312667209043242744224019824380593567642582998924478621582395884770188051376858532702102204361012885895484879752302048075219707736950847555361068281008017371, exp=65537, mod=100753218594801373101605241782117089415967523849664043595259867223687534395978541784644211629212268515702620352659999800812530639439086042593164789038129682257983055916965867275106415277800663102399392424156006808774300993702239063475527499129232811232968510963100403483770572026134850128814034740695252631853";
	REPORT "Expected output is 85923654077259944362850857624610944630400326089823878636524635381935390549840336605379660471462899314317149751023285809596138142553535016420474420073293817183542981215871277711376176316463817598111121213219143738155251327738760275117237355922359111349714288216173788759937613460045194419940190995834815348840, 0111101001011011111111100000100000101011101010011100010111111000110101010111010110110001110111010010111010011000100000111100111110010011011101101001001101100011101011110101101111100111111000100101110010111001010011101100000100101110010010100001100111111010000011100101010010011011101101111100010101001000101000110001001011010101001111010101100001100001001001100101000010101001010001110110011101110111010100010010110110011011010010000100110101011110001111010100100011101101101001011000000111100110010011100100000000010101101010101100110100111101001011100011101101111011100111110010111011101001001001110001101010101110111110101100101010101100110000101000010010010011110010111110001001010111001011101001000101111111001111001110001111101011111111100000010100101110011010111010010101111010110001111011101110000110101011110011011110000010101000101101010010100100111011010010000010001011100001111011110100010001110100100101001110111010011010010111111111000100010011001101111100000001110000011110111011110100110011111000000001101000";
	N_in <= "0100110011111000110010110101100001000101011000110100010101010110011100010001100001011011011000011110101001100011011011001010100011101110001010110000011101010001111110110111001101100011100001011111000001101000001000001001011100010100110101001011100010100001010011000100010101111011100011101011101101101100000111001101101101111101101101010000100010101100011110010100100111101111010101100010110101010010000011010101100101000101001001001110001100000000011001010010110011000111010111000001011111101011100000010000000111100101000011010100001010010010110111110000100011010101110000111111101000110011000011100100011100111001000110101110110000111100010011111010011001001000001110101110011010110110011101110100011110011110110001010111001000001010010010011010001010010000001100101000011101101001100110101011111010010010100010110001011000110101001010001010001100100000100000110111011100110101010001000111001010100000000110010011101110000001001111000011011100001110011101000000001000011111101100001111001011110100010100001100111111011011";
	Exp_in <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "1000111101111010001100110101011000001110110001110111100110111110010101111100111100010101100001110011110001010010110001100111110011100000110001001000110100001101110001011000000101100111100010111001110011011000111100000111010110001011001011110011000011001110110001000010101001111001000000100011111011100001111111000101001111110010010001100001000101100001100111100100110101010111010101111011000101011011101010010011001100101101001111000111000100001100001001100101101110011010001110001000100101001101111001001111010001100010101001101110100010111111000111100100001001001101010101011101101001100001010101000110011101100111101100110110101001101111110011110010111100110100011000111100111110011011010010010101101010111001011110000000001101100001111111100100110011011011000110110010101011110101000011111100001100111101001100010101011101111000111101001110010110100111110110001001001010010010010011011000001110001011110001001001101000011101010011101110000110111011111101111010000001101000011011010100110010000001110000001000000100101101";
	wait for 2102273 * clk_period;
	ASSERT(C_out = "0111101001011011111111100000100000101011101010011100010111111000110101010111010110110001110111010010111010011000100000111100111110010011011101101001001101100011101011110101101111100111111000100101110010111001010011101100000100101110010010100001100111111010000011100101010010011011101101111100010101001000101000110001001011010101001111010101100001100001001001100101000010101001010001110110011101110111010100010010110110011011010010000100110101011110001111010100100011101101101001011000000111100110010011100100000000010101101010101100110100111101001011100011101101111011100111110010111011101001001001110001101010101110111110101100101010101100110000101000010010010011110010111110001001010111001011101001000101111111001111001110001111101011111111100000010100101110011010111010010101111010110001111011101110000110101011110011011110000010101000101101010010100100111011010010000010001011100001111011110100010001110100100101001110111010011010010111111111000100010011001101111100000001110000011110111011110100110011111000000001101000") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=85923654077259944362850857624610944630400326089823878636524635381935390549840336605379660471462899314317149751023285809596138142553535016420474420073293817183542981215871277711376176316463817598111121213219143738155251327738760275117237355922359111349714288216173788759937613460045194419940190995834815348840, exp=12867608215793940718379478366667989660980029214362696566707738966725127224229677811579291870798277117909439436528437345816880257749136368410284097067042427746873568214522605685415681035583560000113540283937701093957956728251956582002489115895815583711917259896866846423964143566160255357197952828427132082873, mod=100753218594801373101605241782117089415967523849664043595259867223687534395978541784644211629212268515702620352659999800812530639439086042593164789038129682257983055916965867275106415277800663102399392424156006808774300993702239063475527499129232811232968510963100403483770572026134850128814034740695252631853";
	REPORT "Expected output is 54051473182883694870366764758765700911582559777313054613910121608584026737001907012426262195401178256691273833725480698483655594641432143815158493354852312667209043242744224019824380593567642582998924478621582395884770188051376858532702102204361012885895484879752302048075219707736950847555361068281008017371, 0100110011111000110010110101100001000101011000110100010101010110011100010001100001011011011000011110101001100011011011001010100011101110001010110000011101010001111110110111001101100011100001011111000001101000001000001001011100010100110101001011100010100001010011000100010101111011100011101011101101101100000111001101101101111101101101010000100010101100011110010100100111101111010101100010110101010010000011010101100101000101001001001110001100000000011001010010110011000111010111000001011111101011100000010000000111100101000011010100001010010010110111110000100011010101110000111111101000110011000011100100011100111001000110101110110000111100010011111010011001001000001110101110011010110110011101110100011110011110110001010111001000001010010010011010001010010000001100101000011101101001100110101011111010010010100010110001011000110101001010001010001100100000100000110111011100110101010001000111001010100000000110010011101110000001001111000011011100001110011101000000001000011111101100001111001011110100010100001100111111011011";
	N_in <= "0111101001011011111111100000100000101011101010011100010111111000110101010111010110110001110111010010111010011000100000111100111110010011011101101001001101100011101011110101101111100111111000100101110010111001010011101100000100101110010010100001100111111010000011100101010010011011101101111100010101001000101000110001001011010101001111010101100001100001001001100101000010101001010001110110011101110111010100010010110110011011010010000100110101011110001111010100100011101101101001011000000111100110010011100100000000010101101010101100110100111101001011100011101101111011100111110010111011101001001001110001101010101110111110101100101010101100110000101000010010010011110010111110001001010111001011101001000101111111001111001110001111101011111111100000010100101110011010111010010101111010110001111011101110000110101011110011011110000010101000101101010010100100111011010010000010001011100001111011110100010001110100100101001110111010011010010111111111000100010011001101111100000001110000011110111011110100110011111000000001101000";
	Exp_in <= "0001001001010010111101110000111101111100100111111011100101001010101110000000100000111000101001011010011011101100101000110111000011111011011110111101111011001111111011010111001110010011011101111101111100110110010011011010111110010101011100010001011101111000101100001101000100000011110101110110011110010100100100010001011101011111100011111101011101010100011100100101010101001010010111000110011011001000011000000001100110101011001000110101011100000100110010000011100101010110101111101101100110010111110011111111010111111111110011110101000101001100111101101111101111111111101101111111011110000101101110100010011100100110001011100111101110001101101111100111110110101010000110000110110111111000101011111101110011110101000001010010100111011100101010111010000010110001111000100110011110001111111110000011111111001111111100000011110001011110100100101001111101011101011110011010110001101000101101000111001111110111001001101011000100000000101111010101001011101110100001001001111000011000110100001001101100011111001011100001101010111001";
	M_in <= "1000111101111010001100110101011000001110110001110111100110111110010101111100111100010101100001110011110001010010110001100111110011100000110001001000110100001101110001011000000101100111100010111001110011011000111100000111010110001011001011110011000011001110110001000010101001111001000000100011111011100001111111000101001111110010010001100001000101100001100111100100110101010111010101111011000101011011101010010011001100101101001111000111000100001100001001100101101110011010001110001000100101001101111001001111010001100010101001101110100010111111000111100100001001001101010101011101101001100001010101000110011101100111101100110110101001101111110011110010111100110100011000111100111110011011010010010101101010111001011110000000001101100001111111100100110011011011000110110010101011110101000011111100001100111101001100010101011101111000111101001110010110100111110110001001001010010010010011011000001110001011110001001001101000011101010011101110000110111011111101111010000001101000011011010100110010000001110000001000000100101101";
	wait for 2102273 * clk_period;
	ASSERT(C_out = "0100110011111000110010110101100001000101011000110100010101010110011100010001100001011011011000011110101001100011011011001010100011101110001010110000011101010001111110110111001101100011100001011111000001101000001000001001011100010100110101001011100010100001010011000100010101111011100011101011101101101100000111001101101101111101101101010000100010101100011110010100100111101111010101100010110101010010000011010101100101000101001001001110001100000000011001010010110011000111010111000001011111101011100000010000000111100101000011010100001010010010110111110000100011010101110000111111101000110011000011100100011100111001000110101110110000111100010011111010011001001000001110101110011010110110011101110100011110011110110001010111001000001010010010011010001010010000001100101000011101101001100110101011111010010010100010110001011000110101001010001010001100100000100000110111011100110101010001000111001010100000000110010011101110000001001111000011011100001110011101000000001000011111101100001111001011110100010100001100111111011011") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=53610029322691035592770787051602554232304283070811234942370481243198510284356840895498134427728655445156946761804583095632225871135156127715795286657675771267940186713831805996946700803831743686492117902608784121609757547378587345679468656034891067994385505920130114395901909229467820330657310634898297904928, exp=65537, mod=96576662507270292424674747143366545500518235781561354837538035391356989209844070999132139779793269203607898511467219515296038152718395572132774968878437700159461036175191384290296121609073326622638247935746347732656460650512661739397752775520253505434182985586410604056699378183286817470413222118941558210829";
	REPORT "Expected output is 11388039982470602092109357764259824395683546510722597370775260417612407365996180232131420872704936172957563864245053618346261253584812498664726885404984005961764491393194497099896856430347871258573910186116334157044156384734478282465339909318243184067696196293620516161944404985681794961366286672292434899416, 0001000000110111100101000101011100010101011000010100111110001010000111111010110000010000011011101000100110111100111101001111110001111001100011101100010010111111100111001010001011110010100101101100100111011110100001010001000010101011100011110111010100011010100001110111111100001011101110111110000110111100011100110000000000101011001001000010101001111010111110000100110001101110001011000011110011100010110010000110111101111100110010000111011111100011110110100101100010111110010110101011011010001010001111111010110110101010001001010100011100010101110001000000110001000101010101000000011010110101000101100000100110111100011000000111111000001011000011001100000110000100100101000111011110000110010001001011001011111111011110010101111000111010110101010011000000100011110001101110100011001001110010100110101011111100000100110100000000011101101100000100110011100011010011010100010000010010110110011111110101001010101000001101010100001010000011111101000101111001011110001001011100010010110100100011001100100111000111110111000111011000";
	N_in <= "0100110001010111110111001111111011010000111100110100111011100101011111000101011001000001101011111010110011111100101011110001101100100111010011010101011110011011101000010001110011110010000001100101111101010001000100001010010110100000001010100000100011010000110000111001111001001001110111100110010100101010011011010001110000001000110111110000001110110011001010111110100101000110110111110010000111100111111001100001111101011111100101011000010111101101111001101010010110000100100010110000000101010010010000110001011100000001011011010000111001101000010010000101101110001010000011011100000100100100111000101000111111110101000000000100011111001110101100010110110010010101111100001011111110001100010110011010000001010001111000000010100011011100000001010000111100011110101100010101110100100000001110011110100010010010010100110100111011000101101010010000111001000111100000000110011110011011111011001010011011011110100011110011101011010011100101100100000000110110010101010111100010001001111111010000110100001101110001101101111100100000";
	Exp_in <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "1000100110000111100111001000110100101011110100100111011000110011000101011110001100010110000100111011011100000010100010101111101011010000011001010111010001011001011010000101000000010001001000010010101011011111001110001000011100011101010111010001011100001010010000110100010111010001101110100100101010001110110001011001101100010010110001101110101011100010000011100101101100100110110000111111000011110011000011011111100010100100011000000001011111001101010000001010100111110001000010010001010110100010001111101000011011101101111000111000000001001001010101001010000001011010110100011000001100110000101001010101000000110101111101010110100101011011111110111000010010111001111001110010000010111101001100011110000010101111001100001100000011101011011101101101000111100011111011100100111100101110010001111101011010001110101111010011010110101110011000111011111011111000011111011001011100110111111111011101101111010010000100011001000010101000010100001011101110110010000011011000011100000101000110110110110110101000100010101000000100001101";
	wait for 2102273 * clk_period;
	ASSERT(C_out = "0001000000110111100101000101011100010101011000010100111110001010000111111010110000010000011011101000100110111100111101001111110001111001100011101100010010111111100111001010001011110010100101101100100111011110100001010001000010101011100011110111010100011010100001110111111100001011101110111110000110111100011100110000000000101011001001000010101001111010111110000100110001101110001011000011110011100010110010000110111101111100110010000111011111100011110110100101100010111110010110101011011010001010001111111010110110101010001001010100011100010101110001000000110001000101010101000000011010110101000101100000100110111100011000000111111000001011000011001100000110000100100101000111011110000110010001001011001011111111011110010101111000111010110101010011000000100011110001101110100011001001110010100110101011111100000100110100000000011101101100000100110011100011010011010100010000010010110110011111110101001010101000001101010100001010000011111101000101111001011110001001011100010010110100100011001100100111000111110111000111011000") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=11388039982470602092109357764259824395683546510722597370775260417612407365996180232131420872704936172957563864245053618346261253584812498664726885404984005961764491393194497099896856430347871258573910186116334157044156384734478282465339909318243184067696196293620516161944404985681794961366286672292434899416, exp=68311148926362538346860896571065193451363708102141662951445949137155264839884824682786356892016674354981884178366028775364498597851808064784578396217862753574486207850976267960844694867854691409669583858236123361380966336068879534279622758130797631283274188888624008402679538184492970760147020718049324624513, mod=96576662507270292424674747143366545500518235781561354837538035391356989209844070999132139779793269203607898511467219515296038152718395572132774968878437700159461036175191384290296121609073326622638247935746347732656460650512661739397752775520253505434182985586410604056699378183286817470413222118941558210829";
	REPORT "Expected output is 53610029322691035592770787051602554232304283070811234942370481243198510284356840895498134427728655445156946761804583095632225871135156127715795286657675771267940186713831805996946700803831743686492117902608784121609757547378587345679468656034891067994385505920130114395901909229467820330657310634898297904928, 0100110001010111110111001111111011010000111100110100111011100101011111000101011001000001101011111010110011111100101011110001101100100111010011010101011110011011101000010001110011110010000001100101111101010001000100001010010110100000001010100000100011010000110000111001111001001001110111100110010100101010011011010001110000001000110111110000001110110011001010111110100101000110110111110010000111100111111001100001111101011111100101011000010111101101111001101010010110000100100010110000000101010010010000110001011100000001011011010000111001101000010010000101101110001010000011011100000100100100111000101000111111110101000000000100011111001110101100010110110010010101111100001011111110001100010110011010000001010001111000000010100011011100000001010000111100011110101100010101110100100000001110011110100010010010010100110100111011000101101010010000111001000111100000000110011110011011111011001010011011011110100011110011101011010011100101100100000000110110010101010111100010001001111111010000110100001101110001101101111100100000";
	N_in <= "0001000000110111100101000101011100010101011000010100111110001010000111111010110000010000011011101000100110111100111101001111110001111001100011101100010010111111100111001010001011110010100101101100100111011110100001010001000010101011100011110111010100011010100001110111111100001011101110111110000110111100011100110000000000101011001001000010101001111010111110000100110001101110001011000011110011100010110010000110111101111100110010000111011111100011110110100101100010111110010110101011011010001010001111111010110110101010001001010100011100010101110001000000110001000101010101000000011010110101000101100000100110111100011000000111111000001011000011001100000110000100100101000111011110000110010001001011001011111111011110010101111000111010110101010011000000100011110001101110100011001001110010100110101011111100000100110100000000011101101100000100110011100011010011010100010000010010110110011111110101001010101000001101010100001010000011111101000101111001011110001001011100010010110100100011001100100111000111110111000111011000";
	Exp_in <= "0110000101000111001111110000000011001100000000100110111000000000111011000111011001010111111000110101001000001011110001100110101001101010100001011001100010101010101101010001001000001101010010111011110010011011011011111100110010000010100001001001101000001011011101000101001000101010011010101110111011011001110101100000010000111110010111111101110100111100010100001001001101000000111101000100111110110110010111000010011110000111011111010100000011011000101110011110100001111010110010010011011101111000101010011100100000000010001101101001111111000101100011111110010110000001001000110000101100011110010000101101010000010000000100011101101111111010000111010011101001111000111100111000111110101111011100000110001100000001101100101100011110111110000111001111010110000010011001011010011110001110101011100001100110110010100111010010011110000010101001010100011000000001110110101000001001100011110110110010101010101011100001010111111111011001011000001001001011011011011111100111011111111111100001001100111010110101110110101110101010000001";
	M_in <= "1000100110000111100111001000110100101011110100100111011000110011000101011110001100010110000100111011011100000010100010101111101011010000011001010111010001011001011010000101000000010001001000010010101011011111001110001000011100011101010111010001011100001010010000110100010111010001101110100100101010001110110001011001101100010010110001101110101011100010000011100101101100100110110000111111000011110011000011011111100010100100011000000001011111001101010000001010100111110001000010010001010110100010001111101000011011101101111000111000000001001001010101001010000001011010110100011000001100110000101001010101000000110101111101010110100101011011111110111000010010111001111001110010000010111101001100011110000010101111001100001100000011101011011101101101000111100011111011100100111100101110010001111101011010001110101111010011010110101110011000111011111011111000011111011001011100110111111111011101101111010010000100011001000010101000010100001011101110110010000011011000011100000101000110110110110110101000100010101000000100001101";
	wait for 2102273 * clk_period;
	ASSERT(C_out = "0100110001010111110111001111111011010000111100110100111011100101011111000101011001000001101011111010110011111100101011110001101100100111010011010101011110011011101000010001110011110010000001100101111101010001000100001010010110100000001010100000100011010000110000111001111001001001110111100110010100101010011011010001110000001000110111110000001110110011001010111110100101000110110111110010000111100111111001100001111101011111100101011000010111101101111001101010010110000100100010110000000101010010010000110001011100000001011011010000111001101000010010000101101110001010000011011100000100100100111000101000111111110101000000000100011111001110101100010110110010010101111100001011111110001100010110011010000001010001111000000010100011011100000001010000111100011110101100010101110100100000001110011110100010010010010100110100111011000101101010010000111001000111100000000110011110011011111011001010011011011110100011110011101011010011100101100100000000110110010101010111100010001001111111010000110100001101110001101101111100100000") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=84398425293680322404764008159378442695079151471103390246281210693416232270315410151342351193652255261082752143396729127398787552054192322636527690462930873820352474641724986444465563912150517736912417041919717808984865461225698798554979308740843650546537837375497770389645958405419532313821141199925014083236, exp=65537, mod=126659643222211502696226346485046946042468021413401959695031378452732557993569430054803022694778819962355629897360446810909544930425107853340851512907898411427721529803299921130934910979359931293511463428232199833579061294764293101259054589379835286815090576263534380922331615656353904133980306913335698449233";
	REPORT "Expected output is 89811918028678530009398645930026705224835015162022731875761285876323316339559183720623980280401285046046868569656377869948211047966888147266835626887568870938051685571049680131184394338792721203273905155733576474872353295339440868108092405447707833278827425959600334040569585206830257062199036461261836032299, 0111111111100101011110111000111101110111011010101001110011111000101110110001010100011001000111111101101100001000111110111000110001000110110101111111111010111001101100110101110110010101111000001000111100110011101110000111010011111000011110110001111111000011110011000010111100101011011000101011101100100000010011001000111111000010010010000100101000000000100111100110110000101010010011011000101001100110010011010001101101010111000111100101110110100100000101101000010011010011100011110010101110101010010011010011001100011110111001111111100010010100001111001111100101011101011010011110001001001101011101111000010001010110001111100110110011110010111100010010111111110011011001010010100100000000111110100111101101010000001100010000100010010110001011101101100000011001111110110001001111000000000001001101010111101110001101111110011101111110101001000101100001010000111010001111110110110101101111010110010010001111111110000001111000101101000000011000010111101000010011010000001101010011001001111101011001101010010010001001100100101011";
	N_in <= "0111100000101111111101011111101010000010100110101100101110110000101110001110110000010011110000011100000101101011001000000010111100001101001011110001100110010101011101110110010111010111110010100111000110001100100101011111001111011011001010101111000111100110001010101111110001011111011010011110101010000000100000011001111010010010001101101101110110010001000101111010101000110111010110011110110001001100110000111000011100101001010010101001001100001100101010111011001110000010100011010110100101000100011001111111010001000001111110011111110101001111011100100100100010100100010110101110100010110001111100101011010010010001000000000000000010001001111100001010001000001001010011111110001100000111111000111001100110011000010010011111110101010111110001111110010011000011100111011000101101001101010000000001110011011111011001111101101001010000010100110101101011101010100011101011110111001010000101000101101010000110100010100010111110111100101010011110010101111011010010110110011111100011011110011111111111111110000110101011011010100100";
	Exp_in <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "1011010001011110100010111011000111110111111001000101011001011011101110011111001101111001001111111101010110101010010100110101100101000110111001101100100010111111110110111101100010110000000101111101001100110110100010001011110101010000011100111000101011110001110011111100000110010100101011001001101110111010010100101001101101111100111011100111011100111010000101000111100001101110011101110001101111110101110110101011001001010011000001100100001111010010100101110100010011011111101110010010000111001011101101011000010100011100101101110000101010001001101000101000000001101000101111110001101001110100101000010011000110101111111001110110101010010010011100001011011011001011100011000100000000011101111110101001110101111010110001110110100100001001100000001110110001111000001110000110110111100100110000011111011110111110110010101110011111100011000001000101010110100111011101100000110111000011101101110110100000001000100011000100110100011010010001101110100111111110010100101100100011011100010010101010110101100011000100101110001101010001";
	wait for 2102273 * clk_period;
	ASSERT(C_out = "0111111111100101011110111000111101110111011010101001110011111000101110110001010100011001000111111101101100001000111110111000110001000110110101111111111010111001101100110101110110010101111000001000111100110011101110000111010011111000011110110001111111000011110011000010111100101011011000101011101100100000010011001000111111000010010010000100101000000000100111100110110000101010010011011000101001100110010011010001101101010111000111100101110110100100000101101000010011010011100011110010101110101010010011010011001100011110111001111111100010010100001111001111100101011101011010011110001001001101011101111000010001010110001111100110110011110010111100010010111111110011011001010010100100000000111110100111101101010000001100010000100010010110001011101101100000011001111110110001001111000000000001001101010111101110001101111110011101111110101001000101100001010000111010001111110110110101101111010110010010001111111110000001111000101101000000011000010111101000010011010000001101010011001001111101011001101010010010001001100100101011") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=89811918028678530009398645930026705224835015162022731875761285876323316339559183720623980280401285046046868569656377869948211047966888147266835626887568870938051685571049680131184394338792721203273905155733576474872353295339440868108092405447707833278827425959600334040569585206830257062199036461261836032299, exp=82199184361919215598454292517234794224304589571613167367274586696852482667538871158137878774651460558751692186009956570511386926176674050052536651841227141433638605108739169310253988214617986946836823227584950059179541616262313659032121088582839764474896488309880083273272989714509038593063989777860973886913, mod=126659643222211502696226346485046946042468021413401959695031378452732557993569430054803022694778819962355629897360446810909544930425107853340851512907898411427721529803299921130934910979359931293511463428232199833579061294764293101259054589379835286815090576263534380922331615656353904133980306913335698449233";
	REPORT "Expected output is 84398425293680322404764008159378442695079151471103390246281210693416232270315410151342351193652255261082752143396729127398787552054192322636527690462930873820352474641724986444465563912150517736912417041919717808984865461225698798554979308740843650546537837375497770389645958405419532313821141199925014083236, 0111100000101111111101011111101010000010100110101100101110110000101110001110110000010011110000011100000101101011001000000010111100001101001011110001100110010101011101110110010111010111110010100111000110001100100101011111001111011011001010101111000111100110001010101111110001011111011010011110101010000000100000011001111010010010001101101101110110010001000101111010101000110111010110011110110001001100110000111000011100101001010010101001001100001100101010111011001110000010100011010110100101000100011001111111010001000001111110011111110101001111011100100100100010100100010110101110100010110001111100101011010010010001000000000000000010001001111100001010001000001001010011111110001100000111111000111001100110011000010010011111110101010111110001111110010011000011100111011000101101001101010000000001110011011111011001111101101001010000010100110101101011101010100011101011110111001010000101000101101010000110100010100010111110111100101010011110010101111011010010110110011111100011011110011111111111111110000110101011011010100100";
	N_in <= "0111111111100101011110111000111101110111011010101001110011111000101110110001010100011001000111111101101100001000111110111000110001000110110101111111111010111001101100110101110110010101111000001000111100110011101110000111010011111000011110110001111111000011110011000010111100101011011000101011101100100000010011001000111111000010010010000100101000000000100111100110110000101010010011011000101001100110010011010001101101010111000111100101110110100100000101101000010011010011100011110010101110101010010011010011001100011110111001111111100010010100001111001111100101011101011010011110001001001101011101111000010001010110001111100110110011110010111100010010111111110011011001010010100100000000111110100111101101010000001100010000100010010110001011101101100000011001111110110001001111000000000001001101010111101110001101111110011101111110101001000101100001010000111010001111110110110101101111010110010010001111111110000001111000101101000000011000010111101000010011010000001101010011001001111101011001101010010010001001100100101011";
	Exp_in <= "0111010100001110001101101101001011010100111100100001011100101001100010000101000001111110100010111111001011111010100010110000010100010001100000101000110100011110000101100110101101010110001111001110000000010010001100000100001111001100100001100110111111010001111001101110011011010110101110011111111010000110101110010011110110110111101000100111101100110101111100100011101100000110010101011011111010001011100110111101011011000111000100101111010111001001001000011110101011001100110101100010110111000100000001010110010111110010100101111000011101010011100110110011011100100011100111110011011100101110101011101110100111011100011000000100100000000001101111110111010000111000100000001010101110110111011001101101000100110111001000101011100110111000101100110010000101010000111101001100111010111001001001100011000010011011010000011100110100000010110110001110010100000001011010110110001110001100010111010001001110010101101111110011010110000111111100001010111111000011111000001101100101011100101110000001111100000010001000001111110111000001";
	M_in <= "1011010001011110100010111011000111110111111001000101011001011011101110011111001101111001001111111101010110101010010100110101100101000110111001101100100010111111110110111101100010110000000101111101001100110110100010001011110101010000011100111000101011110001110011111100000110010100101011001001101110111010010100101001101101111100111011100111011100111010000101000111100001101110011101110001101111110101110110101011001001010011000001100100001111010010100101110100010011011111101110010010000111001011101101011000010100011100101101110000101010001001101000101000000001101000101111110001101001110100101000010011000110101111111001110110101010010010011100001011011011001011100011000100000000011101111110101001110101111010110001110110100100001001100000001110110001111000001110000110110111100100110000011111011110111110110010101110011111100011000001000101010110100111011101100000110111000011101101110110100000001000100011000100110100011010010001101110100111111110010100101100100011011100010010101010110101100011000100101110001101010001";
	wait for 2102273 * clk_period;
	ASSERT(C_out = "0111100000101111111101011111101010000010100110101100101110110000101110001110110000010011110000011100000101101011001000000010111100001101001011110001100110010101011101110110010111010111110010100111000110001100100101011111001111011011001010101111000111100110001010101111110001011111011010011110101010000000100000011001111010010010001101101101110110010001000101111010101000110111010110011110110001001100110000111000011100101001010010101001001100001100101010111011001110000010100011010110100101000100011001111111010001000001111110011111110101001111011100100100100010100100010110101110100010110001111100101011010010010001000000000000000010001001111100001010001000001001010011111110001100000111111000111001100110011000010010011111110101010111110001111110010011000011100111011000101101001101010000000001110011011111011001111101101001010000010100110101101011101010100011101011110111001010000101000101101010000110100010100010111110111100101010011110010101111011010010110110011111100011011110011111111111111110000110101011011010100100") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=53286381971825856799249203420607070528565497649430599643312111847245683787931421411506529846837106464746215507187302760926178478020547521650594973199748292874668820807113680822371833539452016780771592555528849676616990137568792108175600391450928177568007151172437923520993933189629236953777364007808567914192, exp=65537, mod=112929778503919991935446241438216123898434144927734957929381520683898656794503426080108882874737071773575935147348434363190574935911157816005637107284596294482542466331774544931118905224043724185208444257801877481240249742250738950411931346446422038223023266693179946789982520902951606599648238080191667844339";
	REPORT "Expected output is 101393909963639714167179618494089309782974999413426938035232591460151025208952154343665426128144227781779774534433714858570445520940924691293118779975530969554603607703494071785745291033968003680511121915085183182868964237027234412765512266377260032956827729437675415581512854166765659920346706686563530859307, 1001000001100011110001001011101100001110001101100001101000011111100111101001000001111000101001100111010001000100110000010100110011111000110110110000110010100000010110001111000010011011111111011100110110011101000001010000011000101101010000100101110000011100010111011101110001101110100100000101100011011001100110101010101100010100110001010010101000100000000100010011111110011000111001111000100101011001010011011010100111001100111001101001101010111111111100001111011010010101101000011101101000011110001110001001111011110110100001010100111110000011011110011000010001110111000010101101101100010010111001000111101110111000001001110101111011001101110001110110101010110010000010101111000110011111100001111000011010000101010011100101001011010001110100110010110110001000100001001101110101000001110110010100111001111111010001111001011100111001000110010100001110010110111011100001001111111101011101110011111100010010101001011101110100101100100101000100101001111101000111011011111110101011101110010000111111111001111101000110001100101011";
	N_in <= "0100101111100001111000000010101001100100100100100010000000011001101110111001110101101011111010111100010011011110101001000111110111000010011010000101100111001001101100101000111100000101001010000100000010110111111000001101111000001110001000001100011001010010001010011010110011101110010011010100010000010101100010110100011100011100010000101000011110001111110101011100001000011100000000001101000011010010101010101011010010001011000101111011001000010100110011100000110010101000111111000101011001011001100110010100000101111010100010010101000101101010001101111010100101001011110001000100111101011000010110001010110110111110101011000011110100001001000100111010000000110000110110100011010111101000111101101110110001010101011001110000010011111101111100011100011011111111000101111010010001111110010000000101001000011010100111101011000010101010001010011111000000010100001111000011000010000000111100101001001001110011111010111100110110010010101001000011110110111000000110010011100011110111111100110011011011100001010011001010111011010000";
	Exp_in <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "1010000011010001001111010101111101010001010000000011011110000111001011001101111000000011100011100111100111101100010111001110111001101000011111110011000111110100110000101000000011011101100011100010100101001010100011001100000111110010111100100000100010110111100100011110011011011011001111100001101000101011010011001010111101000000011010100000110011001111100111111111000101100111110100110001010111001011110111101101011111110010110000101001000000100011000000001000000110000001011101010011100110001111100001100011011101111000101001101111100100010011100010100101000010011001000100111111000101010001100010110001001001010001110110011000001011000011101000001011001101101101101110010011100101110101110111110000011110100001100011011001100110101110010010110000000011001110001100011101110101010011000011000110010000010011011010000001111100100110100111110001011001011111000000000001010010000110110110011110000011011001110001101111001100111100001001110000010100011001011101000100111001100101101111011011101001010111111010110011010011110011";
	wait for 2102273 * clk_period;
	ASSERT(C_out = "1001000001100011110001001011101100001110001101100001101000011111100111101001000001111000101001100111010001000100110000010100110011111000110110110000110010100000010110001111000010011011111111011100110110011101000001010000011000101101010000100101110000011100010111011101110001101110100100000101100011011001100110101010101100010100110001010010101000100000000100010011111110011000111001111000100101011001010011011010100111001100111001101001101010111111111100001111011010010101101000011101101000011110001110001001111011110110100001010100111110000011011110011000010001110111000010101101101100010010111001000111101110111000001001110101111011001101110001110110101010110010000010101111000110011111100001111000011010000101010011100101001011010001110100110010110110001000100001001101110101000001110110010100111001111111010001111001011100111001000110010100001110010110111011100001001111111101011101110011111100010010101001011101110100101100100101000100101001111101000111011011111110101011101110010000111111111001111101000110001100101011") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=101393909963639714167179618494089309782974999413426938035232591460151025208952154343665426128144227781779774534433714858570445520940924691293118779975530969554603607703494071785745291033968003680511121915085183182868964237027234412765512266377260032956827729437675415581512854166765659920346706686563530859307, exp=93608149403343907134918925490786162239018210919850982720535296544426974559479440901717120913182121351720998839503736032256050670894879796095186351050122742617457290010720110668232518831932496084397709562823876246343346622946920137924933293844041763590192372926226569621397916402691663075923231258885577914593, mod=112929778503919991935446241438216123898434144927734957929381520683898656794503426080108882874737071773575935147348434363190574935911157816005637107284596294482542466331774544931118905224043724185208444257801877481240249742250738950411931346446422038223023266693179946789982520902951606599648238080191667844339";
	REPORT "Expected output is 53286381971825856799249203420607070528565497649430599643312111847245683787931421411506529846837106464746215507187302760926178478020547521650594973199748292874668820807113680822371833539452016780771592555528849676616990137568792108175600391450928177568007151172437923520993933189629236953777364007808567914192, 0100101111100001111000000010101001100100100100100010000000011001101110111001110101101011111010111100010011011110101001000111110111000010011010000101100111001001101100101000111100000101001010000100000010110111111000001101111000001110001000001100011001010010001010011010110011101110010011010100010000010101100010110100011100011100010000101000011110001111110101011100001000011100000000001101000011010010101010101011010010001011000101111011001000010100110011100000110010101000111111000101011001011001100110010100000101111010100010010101000101101010001101111010100101001011110001000100111101011000010110001010110110111110101011000011110100001001000100111010000000110000110110100011010111101000111101101110110001010101011001110000010011111101111100011100011011111111000101111010010001111110010000000101001000011010100111101011000010101010001010011111000000010100001111000011000010000000111100101001001001110011111010111100110110010010101001000011110110111000000110010011100011110111111100110011011011100001010011001010111011010000";
	N_in <= "1001000001100011110001001011101100001110001101100001101000011111100111101001000001111000101001100111010001000100110000010100110011111000110110110000110010100000010110001111000010011011111111011100110110011101000001010000011000101101010000100101110000011100010111011101110001101110100100000101100011011001100110101010101100010100110001010010101000100000000100010011111110011000111001111000100101011001010011011010100111001100111001101001101010111111111100001111011010010101101000011101101000011110001110001001111011110110100001010100111110000011011110011000010001110111000010101101101100010010111001000111101110111000001001110101111011001101110001110110101010110010000010101111000110011111100001111000011010000101010011100101001011010001110100110010110110001000100001001101110101000001110110010100111001111111010001111001011100111001000110010100001110010110111011100001001111111101011101110011111100010010101001011101110100101100100101000100101001111101000111011011111110101011101110010000111111111001111101000110001100101011";
	Exp_in <= "1000010101001101011011000000010111111010100111111011010001100111100001000011010101110011110101010100001000010011001111101110010100010000000100010111111100100011010101111010011011100001111111111101100100010010010001101010001011101101111100101101101001101110111011111010110111100000110001100001010110000011000101101100100110011110001001110100100111111111010000001010000100100110011000101011111010001010100000110110100110010101011111001101100101100101011010100010000111101111011000001101001000111010011110011111010110110000100111010100111110000010110110111101000110100110110100101101100010101000111000000010011010101000100110010010011101001001010011011010100111110111100011100101110000101011001101000111111111011101001001001001101000110110101111111010100111110100111001011111111010101001000100000000100101100000000110010111111000010010111101100111101111111010010111100001000101010010011000001010100111011110101011000100101011101101011000010000101011110011111010001111000110000111111110010011001010011011011100100011100011100001";
	M_in <= "1010000011010001001111010101111101010001010000000011011110000111001011001101111000000011100011100111100111101100010111001110111001101000011111110011000111110100110000101000000011011101100011100010100101001010100011001100000111110010111100100000100010110111100100011110011011011011001111100001101000101011010011001010111101000000011010100000110011001111100111111111000101100111110100110001010111001011110111101101011111110010110000101001000000100011000000001000000110000001011101010011100110001111100001100011011101111000101001101111100100010011100010100101000010011001000100111111000101010001100010110001001001010001110110011000001011000011101000001011001101101101101110010011100101110101110111110000011110100001100011011001100110101110010010110000000011001110001100011101110101010011000011000110010000010011011010000001111100100110100111110001011001011111000000000001010010000110110110011110000011011001110001101111001100111100001001110000010100011001011101000100111001100101101111011011101001010111111010110011010011110011";
	wait for 2102273 * clk_period;
	ASSERT(C_out = "0100101111100001111000000010101001100100100100100010000000011001101110111001110101101011111010111100010011011110101001000111110111000010011010000101100111001001101100101000111100000101001010000100000010110111111000001101111000001110001000001100011001010010001010011010110011101110010011010100010000010101100010110100011100011100010000101000011110001111110101011100001000011100000000001101000011010010101010101011010010001011000101111011001000010100110011100000110010101000111111000101011001011001100110010100000101111010100010010101000101101010001101111010100101001011110001000100111101011000010110001010110110111110101011000011110100001001000100111010000000110000110110100011010111101000111101101110110001010101011001110000010011111101111100011100011011111111000101111010010001111110010000000101001000011010100111101011000010101010001010011111000000010100001111000011000010000000111100101001001001110011111010111100110110010010101001000011110110111000000110010011100011110111111100110011011011100001010011001010111011010000") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=64828386337539654265576501996577739565702775771988394226504455907473226577420635153447751505878294031955541862866357208477685703915994468171609280166427890237321754467345968101738171539531597457506866748878785388802038810027406685305610061890576890717635490763593633374657679905292609842840054378702565435835, exp=65537, mod=108015386519967823516896221166170740556607682492638988243544873291461732283801943917361169164582973418809395231987761972573718992936095557711738159719491681765007268734766305990898363604648973311687835858810239324522834597975978924037258740009701811170349169459266226425901140999993463829165833856884308205503";
	REPORT "Expected output is 2068257946745193880534535393793905638057274071566901597119644136973453745791060699260005141085689930702317674047099482404121088276135240280816390493062997168020104380352258984632389035626239918944881322204164549784207253343675856736696381886811340222747169365860874285925430656948222428647697271802251607766, 0000001011110001111111101111110101010010010110001000000000011101100010001001100011001110100110111110100000110101101101110011011001001111111100010001011110001000011111010101101110100001101101011101111000101110100011001011100111110011111110001010100001110100000010100101100000111111000011110001001000110100000110101110110100110011000100001011001110001111100010010111101110111000001011101100101010101000001101100000100000011011011111000011111000100111100001011111001111011110101110001010110100111011100100111011100000101110011011001111110101111111111101010000010010000100011011101000111100111110100011000010110001010010110011110101000111100010010001001101110100010000000010100010000010010000000010011010110011000011000000010100101011001001001010111101001000000001010100010000010000011100110011000110011011011101000110011001111111010000000001011010001010100100000100001011111010001011101101000110101101110111110101101010111001000011011110111101101001000000100110110100010001111100100101111101101110000100010101100111111011010110";
	N_in <= "0101110001010001100101010111000100000110110001110110110100110101011001001111100111101110100111001000011011010011000111101000000000111100100010111101110011011000101001000000111001011110000000110100110011101011110100101001010001101111001000010001001001100010110001101111010101011100000110110011011001010111110100100010010110101010111011011110010001011010100000100100111101100010111000110001100000000000010111110100010111010010011100000101110001100001110101011011111010011100000110001111000100010100001100110111110000110001111001101001100110101101001001101000101010100101110110010010111110110100101011110111100110111000001011011011000111010011111111101010110110110111101111011111101111101101010100000110010001011011100000010101011001100000011000000100101000110100001100001011111111011101011111111111011100100100100010011011101101000111011101001111001001011011001010101001110001111100000000100110100000011011011100011101110001001001101010100100001100100011100000101101000000001111100001011110011010101101001000100110100110111011";
	Exp_in <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "1001100111010001101010110000110000111010010100100000001110100011100010001101101001011110010001100010000111110010101100000000110110011010001001000100110001100010001111011001110011111010111011010111010010100110100000011011000010100101101000110100111001000001100001100111000011010000010010110010011100101001101100000001110101001101010000111000001010100101111100000000000111111001000100000111000001100000100111010110001010100011100000110001010001001011001100100101110000110101011011101111011000110101000111110000011111101011111101010011111110000110101101110001110001100000111100011001110010011010011010000001010001000111010001101010000011100001001111111010000101001011111110101110111101001010000000111000111111011011111010100101101111011010000001011011101100000101001111111100001001111110101001101010111110001010110011100111000010100010011100011101011000011111111000001001001110010010001011100101010101010000011001001101111000000001000101110111001110000100000011000100111111111100001010100110010110111101010010000101111110111111";
	wait for 2102273 * clk_period;
	ASSERT(C_out = "0000001011110001111111101111110101010010010110001000000000011101100010001001100011001110100110111110100000110101101101110011011001001111111100010001011110001000011111010101101110100001101101011101111000101110100011001011100111110011111110001010100001110100000010100101100000111111000011110001001000110100000110101110110100110011000100001011001110001111100010010111101110111000001011101100101010101000001101100000100000011011011111000011111000100111100001011111001111011110101110001010110100111011100100111011100000101110011011001111110101111111111101010000010010000100011011101000111100111110100011000010110001010010110011110101000111100010010001001101110100010000000010100010000010010000000010011010110011000011000000010100101011001001001010111101001000000001010100010000010000011100110011000110011011011101000110011001111111010000000001011010001010100100000100001011111010001011101101000110101101110111110101101010111001000011011110111101101001000000100110110100010001111100100101111101101110000100010101100111111011010110") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=2068257946745193880534535393793905638057274071566901597119644136973453745791060699260005141085689930702317674047099482404121088276135240280816390493062997168020104380352258984632389035626239918944881322204164549784207253343675856736696381886811340222747169365860874285925430656948222428647697271802251607766, exp=15545434268525207309021852663980994322747816672575353420405499868548561253960662450654600417479387297041521824741879715661615843590235337295529455388420759466912760551851165769873011463344011308948695220550245316311907540697248635838844306379011901664742124315355593494001025724840870995416040143310309069633, mod=108015386519967823516896221166170740556607682492638988243544873291461732283801943917361169164582973418809395231987761972573718992936095557711738159719491681765007268734766305990898363604648973311687835858810239324522834597975978924037258740009701811170349169459266226425901140999993463829165833856884308205503";
	REPORT "Expected output is 64828386337539654265576501996577739565702775771988394226504455907473226577420635153447751505878294031955541862866357208477685703915994468171609280166427890237321754467345968101738171539531597457506866748878785388802038810027406685305610061890576890717635490763593633374657679905292609842840054378702565435835, 0101110001010001100101010111000100000110110001110110110100110101011001001111100111101110100111001000011011010011000111101000000000111100100010111101110011011000101001000000111001011110000000110100110011101011110100101001010001101111001000010001001001100010110001101111010101011100000110110011011001010111110100100010010110101010111011011110010001011010100000100100111101100010111000110001100000000000010111110100010111010010011100000101110001100001110101011011111010011100000110001111000100010100001100110111110000110001111001101001100110101101001001101000101010100101110110010010111110110100101011110111100110111000001011011011000111010011111111101010110110110111101111011111101111101101010100000110010001011011100000010101011001100000011000000100101000110100001100001011111111011101011111111111011100100100100010011011101101000111011101001111001001011011001010101001110001111100000000100110100000011011011100011101110001001001101010100100001100100011100000101101000000001111100001011110011010101101001000100110100110111011";
	N_in <= "0000001011110001111111101111110101010010010110001000000000011101100010001001100011001110100110111110100000110101101101110011011001001111111100010001011110001000011111010101101110100001101101011101111000101110100011001011100111110011111110001010100001110100000010100101100000111111000011110001001000110100000110101110110100110011000100001011001110001111100010010111101110111000001011101100101010101000001101100000100000011011011111000011111000100111100001011111001111011110101110001010110100111011100100111011100000101110011011001111110101111111111101010000010010000100011011101000111100111110100011000010110001010010110011110101000111100010010001001101110100010000000010100010000010010000000010011010110011000011000000010100101011001001001010111101001000000001010100010000010000011100110011000110011011011101000110011001111111010000000001011010001010100100000100001011111010001011101101000110101101110111110101101010111001000011011110111101101001000000100110110100010001111100100101111101101110000100010101100111111011010110";
	Exp_in <= "0001011000100011001011101101001011011011101100011110001000000100001011110011010111111110010010110110100110100111010110111101111100011001010010000001000000010110001100110111011111011100010001010100000001111100100101100011110110101110000110010000101010110010001100110111111100011000111110110011011111101111101100000000000100000111100101011010011110111111111010100000001011011110101011011001011011111110110100001010011111011001100100001000101111100011001001101010010001001110101011000100011000011111011111000100111010001011010101011101110010000100111101110101000110100100101001001010111010001001001000110010111110110100101011100010011000110110010101110100001011000011110011111111001110110000101010111011100010110110011110101111110010011011010111011001010101101010101110011000111100110111101101000010000011010101111011110101000100110111000110101000000010100100001101100011001000010100011010011001011000101011101110000001010100101001010111011001011100001010100111111110101110001010011011100001001001110111011101001001001101000001";
	M_in <= "1001100111010001101010110000110000111010010100100000001110100011100010001101101001011110010001100010000111110010101100000000110110011010001001000100110001100010001111011001110011111010111011010111010010100110100000011011000010100101101000110100111001000001100001100111000011010000010010110010011100101001101100000001110101001101010000111000001010100101111100000000000111111001000100000111000001100000100111010110001010100011100000110001010001001011001100100101110000110101011011101111011000110101000111110000011111101011111101010011111110000110101101110001110001100000111100011001110010011010011010000001010001000111010001101010000011100001001111111010000101001011111110101110111101001010000000111000111111011011111010100101101111011010000001011011101100000101001111111100001001111110101001101010111110001010110011100111000010100010011100011101011000011111111000001001001110010010001011100101010101010000011001001101111000000001000101110111001110000100000011000100111111111100001010100110010110111101010010000101111110111111";
	wait for 2102273 * clk_period;
	ASSERT(C_out = "0101110001010001100101010111000100000110110001110110110100110101011001001111100111101110100111001000011011010011000111101000000000111100100010111101110011011000101001000000111001011110000000110100110011101011110100101001010001101111001000010001001001100010110001101111010101011100000110110011011001010111110100100010010110101010111011011110010001011010100000100100111101100010111000110001100000000000010111110100010111010010011100000101110001100001110101011011111010011100000110001111000100010100001100110111110000110001111001101001100110101101001001101000101010100101110110010010111110110100101011110111100110111000001011011011000111010011111111101010110110110111101111011111101111101101010100000110010001011011100000010101011001100000011000000100101000110100001100001011111111011101011111111111011100100100100010011011101101000111011101001111001001011011001010101001110001111100000000100110100000011011011100011101110001001001101010100100001100100011100000101101000000001111100001011110011010101101001000100110100110111011") REPORT "test failed" SEVERITY NOTE;

	wait;

end process;
end;

-- Entity name: modular_exponentiation_tb
-- Author: Luis Gallet, Jacob Barnett
-- Contact: luis.galletzambrano@mail.mcgill.ca, jacob.barnett@mail.mcgill.ca
-- Date: April 06, 2016
-- Description:

library ieee;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
--use IEEE.std_logic_arith.all;
--use IEEE.std_logic_unsigned.all;

entity modular_exponentiation_tb is
end entity;

architecture test of modular_exponentiation_tb is
-- define the ALU compontent to be tested
component modular_exponentiation is
 	generic(
		WIDTH_IN : integer := 64
	);
	port(	N :	in unsigned(WIDTH_IN-1 downto 0); --Number
		Exp :	in unsigned(WIDTH_IN-1 downto 0); --Exponent
		M :	in unsigned(WIDTH_IN-1 downto 0); --Modulus
		--latch_in: in std_logic;
		clk :	in std_logic;
		reset :	in std_logic;
		C : 	out unsigned(WIDTH_IN-1 downto 0) --Output
		--C : out std_logic
	);

end component;

CONSTANT WIDTH_IN : integer := 64;

CONSTANT clk_period : time := 1 ns;

Signal M_in : unsigned(WIDTH_IN-1 downto 0) := (WIDTH_IN-1 downto 0 => '0');
Signal N_in : unsigned(WIDTH_IN-1 downto 0) := (WIDTH_IN-1 downto 0 => '0');
Signal Exp_in : unsigned(WIDTH_IN-1 downto 0) := (WIDTH_IN-1 downto 0 => '0');
signal latch_in : std_logic := '0';

Signal clk : std_logic := '0';
Signal reset_t : std_logic := '0';

Signal C_out : unsigned(WIDTH_IN-1 downto 0) := (WIDTH_IN-1 downto 0 => '0');
--signal c_out : std_logic;

Begin
-- device under test
dut: modular_exponentiation 
			generic map(WIDTH_IN => WIDTH_IN)
			PORT MAP(	N	=> 	N_in,
					Exp 	=> 	Exp_in,
					M 	=> 	M_in,
					--latch_in => latch_in,
					clk	=> 	clk,
					reset 	=>	reset_t,
					C	=>	C_out
				);
  
-- process for clock
clk_process : Process
Begin
	clk <= '0';
	wait for clk_period/2;
	clk <= '1';
	wait for clk_period/2;
end process;

stim_process: process
Begin


	reset_t <= '1';
	wait for 1 * clk_period;
	reset_t <= '0';
	wait for 1 * clk_period;


	REPORT "Begin test case for base=5903434394152496440, exp=65537, mod=10061957843532492581";
	REPORT "Expected output is 3393152870111853512, 0010111100010110111001101000111011000011100111010011101111001000";
	N_in <= "0101000111101101001101100100110111000010010010000110110100111000";
	Exp_in <= "0000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "1000101110100011010000010101100100100000101101011010111100100101";
	wait for 8513 * clk_period;
	ASSERT(C_out = "0010111100010110111001101000111011000011100111010011101111001000") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=3393152870111853512, exp=446775062781666473, mod=10061957843532492581";
	REPORT "Expected output is 5903434394152496440, 0101000111101101001101100100110111000010010010000110110100111000";
	N_in <= "0010111100010110111001101000111011000011100111010011101111001000";
	Exp_in <= "0000011000110011010000111000110101101111100110101010010010101001";
	M_in <= "1000101110100011010000010101100100100000101101011010111100100101";
	wait for 8513 * clk_period;
	ASSERT(C_out = "0101000111101101001101100100110111000010010010000110110100111000") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=6817527486901138695, exp=65537, mod=9541397238521654791";
	REPORT "Expected output is 1638934027748418114, 0001011010111110101010011101000010010110001111101010001001000010";
	N_in <= "0101111010011100101110010010000011100111001101000011010100000111";
	Exp_in <= "0000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "1000010001101001110110100011110001100110111110011110111000000111";
	wait for 8513 * clk_period;
	ASSERT(C_out = "0001011010111110101010011101000010010110001111101010001001000010") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=1638934027748418114, exp=598948810554944497, mod=9541397238521654791";
	REPORT "Expected output is 6817527486901138695, 0101111010011100101110010010000011100111001101000011010100000111";
	N_in <= "0001011010111110101010011101000010010110001111101010001001000010";
	Exp_in <= "0000100001001111111001001100010100010011110001010010101111110001";
	M_in <= "1000010001101001110110100011110001100110111110011110111000000111";
	wait for 8513 * clk_period;
	ASSERT(C_out = "0101111010011100101110010010000011100111001101000011010100000111") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=5228736734326626413, exp=65537, mod=12104320301824256147";
	REPORT "Expected output is 3142956270292174682, 0010101110011110000001100001001101100011010110100000011101011010";
	N_in <= "0100100010010000001101000101101101011001100100110001100001101101";
	Exp_in <= "0000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "1010011111111011001011110010111011011101110010001010100010010011";
	wait for 8513 * clk_period;
	ASSERT(C_out = "0010101110011110000001100001001101100011010110100000011101011010") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=3142956270292174682, exp=3610961226293098193, mod=12104320301824256147";
	REPORT "Expected output is 5228736734326626413, 0100100010010000001101000101101101011001100100110001100001101101";
	N_in <= "0010101110011110000001100001001101100011010110100000011101011010";
	Exp_in <= "0011001000011100101101100001101010000110111010001011011011010001";
	M_in <= "1010011111111011001011110010111011011101110010001010100010010011";
	wait for 8513 * clk_period;
	ASSERT(C_out = "0100100010010000001101000101101101011001100100110001100001101101") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=9118569000187643702, exp=65537, mod=9672413179721907337";
	REPORT "Expected output is 427488509584743641, 0000010111101110101111101000100011010111010111000001110011011001";
	N_in <= "0111111010001011101010100011000110000100000100101100011100110110";
	Exp_in <= "0000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "1000011000111011010100001000101001010010001000010111110010001001";
	wait for 8513 * clk_period;
	ASSERT(C_out = "0000010111101110101111101000100011010111010111000001110011011001") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=427488509584743641, exp=3447190965790685393, mod=9672413179721907337";
	REPORT "Expected output is 9118569000187643702, 0111111010001011101010100011000110000100000100101100011100110110";
	N_in <= "0000010111101110101111101000100011010111010111000001110011011001";
	Exp_in <= "0010111111010110111000011110101101011100111000111011100011010001";
	M_in <= "1000011000111011010100001000101001010010001000010111110010001001";
	wait for 8513 * clk_period;
	ASSERT(C_out = "0111111010001011101010100011000110000100000100101100011100110110") REPORT "test failed" SEVERITY NOTE;




	wait;

end process;
end;

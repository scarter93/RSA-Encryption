-- Entity name: modular_exponentiation_tb
-- Author: Luis Gallet, Jacob Barnett
-- Contact: luis.galletzambrano@mail.mcgill.ca, jacob.barnett@mail.mcgill.ca
-- Date: April 06, 2016
-- Description:

library ieee;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
--use IEEE.std_logic_arith.all;
--use IEEE.std_logic_unsigned.all;

entity modular_exponentiation_tb is
end entity;

architecture test of modular_exponentiation_tb is
-- define the ALU compontent to be tested
component modular_exponentiation is
 	generic(
		WIDTH_IN : integer := 64
	);
	port(	N :	in unsigned(WIDTH_IN-1 downto 0); --Number
		Exp :	in unsigned(WIDTH_IN-1 downto 0); --Exponent
		M :	in unsigned(WIDTH_IN-1 downto 0); --Modulus
		--latch_in: in std_logic;
		clk :	in std_logic;
		reset :	in std_logic;
		C : 	out unsigned(WIDTH_IN-1 downto 0) --Output
		--C : out std_logic
	);

end component;

CONSTANT WIDTH_IN : integer := 64;

CONSTANT clk_period : time := 1 ns;

Signal M_in : unsigned(WIDTH_IN-1 downto 0) := (WIDTH_IN-1 downto 0 => '0');
Signal N_in : unsigned(WIDTH_IN-1 downto 0) := (WIDTH_IN-1 downto 0 => '0');
Signal Exp_in : unsigned(WIDTH_IN-1 downto 0) := (WIDTH_IN-1 downto 0 => '0');
signal latch_in : std_logic := '0';

Signal clk : std_logic := '0';
Signal reset_t : std_logic := '0';

Signal C_out : unsigned(WIDTH_IN-1 downto 0) := (WIDTH_IN-1 downto 0 => '0');
--signal c_out : std_logic;

Begin
-- device under test
dut: modular_exponentiation 
			generic map(WIDTH_IN => WIDTH_IN)
			PORT MAP(	N	=> 	N_in,
					Exp 	=> 	Exp_in,
					M 	=> 	M_in,
					--latch_in => latch_in,
					clk	=> 	clk,
					reset 	=>	reset_t,
					C	=>	C_out
				);
  
-- process for clock
clk_process : Process
Begin
	clk <= '0';
	wait for clk_period/2;
	clk <= '1';
	wait for clk_period/2;
end process;

stim_process: process
Begin


	reset_t <= '1';
	wait for 1 * clk_period;
	reset_t <= '0';
	wait for 1 * clk_period;


	REPORT "Begin test case for base=1475272348399831930, exp=65537, mod=2852210150436973297";
	REPORT "Expected output is 51108437778217609, 0000000010110101100100101101101001110110110010111011101010001001";
	N_in <= "0001010001111001001110000110001001110001010101000000101101111010";
	Exp_in <= "0000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "0010011110010101000101100000010100101001100011110010101011110001";
	wait for 8513 * clk_period;
	ASSERT(C_out = "0000000010110101100100101101101001110110110010111011101010001001") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=51108437778217609, exp=1022647268164012937, mod=2852210150436973297";
	REPORT "Expected output is 1475272348399831930, 0001010001111001001110000110001001110001010101000000101101111010";
	N_in <= "0000000010110101100100101101101001110110110010111011101010001001";
	Exp_in <= "0000111000110001001011000100010110101101011100001000101110001001";
	M_in <= "0010011110010101000101100000010100101001100011110010101011110001";
	wait for 8513 * clk_period;
	ASSERT(C_out = "0001010001111001001110000110001001110001010101000000101101111010") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=2262921332397090273, exp=65537, mod=3097013873315263543";
	REPORT "Expected output is 1136320092719957865, 0000111111000101000001010001101010010101101101100100011101101001";
	N_in <= "0001111101100111100000101111011001011100001011101010010111100001";
	Exp_in <= "0000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "0010101011111010110011011011010110000111011010011011010000110111";
	wait for 8513 * clk_period;
	ASSERT(C_out = "0000111111000101000001010001101010010101101101100100011101101001") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=1136320092719957865, exp=1743036095025014873, mod=3097013873315263543";
	REPORT "Expected output is 2262921332397090273, 0001111101100111100000101111011001011100001011101010010111100001";
	N_in <= "0000111111000101000001010001101010010101101101100100011101101001";
	Exp_in <= "0001100000110000100000100001011111101010101001100110100001011001";
	M_in <= "0010101011111010110011011011010110000111011010011011010000110111";
	wait for 8513 * clk_period;
	ASSERT(C_out = "0001111101100111100000101111011001011100001011101010010111100001") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=1552948844763863111, exp=65537, mod=2579020524292604741";
	REPORT "Expected output is 1313051723566648797, 0001001000111000111001011001010111110010111001111000110111011101";
	N_in <= "0001010110001101001011101011111100010110100000001101100001000111";
	Exp_in <= "0000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "0010001111001010100001011000000010101010111001110000001101000101";
	wait for 8513 * clk_period;
	ASSERT(C_out = "0001001000111000111001011001010111110010111001111000110111011101") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=1313051723566648797, exp=2318037196379765453, mod=2579020524292604741";
	REPORT "Expected output is 1552948844763863111, 0001010110001101001011101011111100010110100000001101100001000111";
	N_in <= "0001001000111000111001011001010111110010111001111000110111011101";
	Exp_in <= "0010000000101011010100101000110001110010010110111011101011001101";
	M_in <= "0010001111001010100001011000000010101010111001110000001101000101";
	wait for 8513 * clk_period;
	ASSERT(C_out = "0001010110001101001011101011111100010110100000001101100001000111") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=2010024926487313335, exp=65537, mod=2516764108772381051";
	REPORT "Expected output is 848932322797645510, 0000101111001000000000110111001100100010101100110110111011000110";
	N_in <= "0001101111100101000010110000010101100100111101001111101110110111";
	Exp_in <= "0000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "0010001011101101010101111001111101011110110101001001000101111011";
	wait for 8513 * clk_period;
	ASSERT(C_out = "0000101111001000000000110111001100100010101100110110111011000110") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=848932322797645510, exp=1045000302219383873, mod=2516764108772381051";
	REPORT "Expected output is 2010024926487313335, 0001101111100101000010110000010101100100111101001111101110110111";
	N_in <= "0000101111001000000000110111001100100010101100110110111011000110";
	Exp_in <= "0000111010000000100101100011110011111011111101100101010001000001";
	M_in <= "0010001011101101010101111001111101011110110101001001000101111011";
	wait for 8513 * clk_period;
	ASSERT(C_out = "0001101111100101000010110000010101100100111101001111101110110111") REPORT "test failed" SEVERITY NOTE;




	wait;

end process;
end;

-- Entity name: modular_exponentiation_tb
-- Author: Luis Gallet, Jacob Barnett
-- Contact: luis.galletzambrano@mail.mcgill.ca, jacob.barnett@mail.mcgill.ca
-- Date: April 09, 2016
-- Description:

library ieee;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
--use IEEE.std_logic_arith.all;
--use IEEE.std_logic_unsigned.all;

entity modular_exponentiation_tb is
end entity;

architecture test of modular_exponentiation_tb is
-- define the ALU compontent to be tested
component modular_exponentiation is
 	generic(
		WIDTH_IN : integer := 128
	);
	port(	N :	in unsigned(WIDTH_IN-1 downto 0); --Number
		Exp :	in unsigned(WIDTH_IN-1 downto 0); --Exponent
		M :	in unsigned(WIDTH_IN-1 downto 0); --Modulus
		--latch_in: in std_logic;
		clk :	in std_logic;
		reset :	in std_logic;
		C : 	out unsigned(WIDTH_IN-1 downto 0) --Output
		--C : out std_logic
	);

end component;

CONSTANT WIDTH_IN : integer := 128;

CONSTANT clk_period : time := 1 ns;

Signal M_in : unsigned(WIDTH_IN-1 downto 0) := (WIDTH_IN-1 downto 0 => '0');
Signal N_in : unsigned(WIDTH_IN-1 downto 0) := (WIDTH_IN-1 downto 0 => '0');
Signal Exp_in : unsigned(WIDTH_IN-1 downto 0) := (WIDTH_IN-1 downto 0 => '0');
signal latch_in : std_logic := '0';

Signal clk : std_logic := '0';
Signal reset_t : std_logic := '0';

Signal C_out : unsigned(WIDTH_IN-1 downto 0) := (WIDTH_IN-1 downto 0 => '0');
--signal c_out : std_logic;

Begin
-- device under test
dut: modular_exponentiation 
			generic map(WIDTH_IN => WIDTH_IN)
			PORT MAP(	N	=> 	N_in,
					Exp 	=> 	Exp_in,
					M 	=> 	M_in,
					--latch_in => latch_in,
					clk	=> 	clk,
					reset 	=>	reset_t,
					C	=>	C_out
				);
  
-- process for clock
clk_process : Process
Begin
	clk <= '0';
	wait for clk_period/2;
	clk <= '1';
	wait for clk_period/2;
end process;

stim_process: process
Begin


	reset_t <= '1';
	wait for 1 * clk_period;
	reset_t <= '0';
	wait for 1 * clk_period;


	REPORT "Begin test case for base=114396660566281941370247871186287366465, exp=65537, mod=192560265107138277498349449196845774883";
	REPORT "Expected output is 136783107359261161669828512609463200599, 01100110111001110111011111011110001111101111010000110010000001011110010100111111010111010110111011010010111100000110101101010111";
	N_in <= "01010110000011111111111011010011010101100101010111100001110011001110110111000001111011011000011011000010010111101001000101000001";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10010000110111011100001000010000101011000001100000001010101010001000111110001110101110011011000011110010101100011011100000100011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01100110111001110111011111011110001111101111010000110010000001011110010100111111010111010110111011010010111100000110101101010111") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=136783107359261161669828512609463200599, exp=11843850476019262333094581869024614817, mod=192560265107138277498349449196845774883";
	REPORT "Expected output is 114396660566281941370247871186287366465, 01010110000011111111111011010011010101100101010111100001110011001110110111000001111011011000011011000010010111101001000101000001";
	N_in <= "01100110111001110111011111011110001111101111010000110010000001011110010100111111010111010110111011010010111100000110101101010111";
	Exp_in <= "00001000111010010000101011101001101110011001110000010100111100101101110001000001110000000011000011011001001110111001100110100001";
	M_in <= "10010000110111011100001000010000101011000001100000001010101010001000111110001110101110011011000011110010101100011011100000100011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01010110000011111111111011010011010101100101010111100001110011001110110111000001111011011000011011000010010111101001000101000001") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=122624919106256087630111067424141196536, exp=65537, mod=179114200985125995187613225846699555213";
	REPORT "Expected output is 66581388608736170524710731800441889647, 00110010000101110001101111100111110100011111010110010000100010100111110100001001010101101001111111100110110110011010001101101111";
	N_in <= "01011100010000001011001101001011000001010110001001100000101000110010001001010010000101000101110101000010100001011011110011111000";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10000110110000000010001111101011101000100000111010100010001110100110011100010010100101101111101001101010100010010111100110001101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "00110010000101110001101111100111110100011111010110010000100010100111110100001001010101101001111111100110110110011010001101101111") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=66581388608736170524710731800441889647, exp=140570361985885384198038659070397650713, mod=179114200985125995187613225846699555213";
	REPORT "Expected output is 122624919106256087630111067424141196536, 01011100010000001011001101001011000001010110001001100000101000110010001001010010000101000101110101000010100001011011110011111000";
	N_in <= "00110010000101110001101111100111110100011111010110010000100010100111110100001001010101101001111111100110110110011010001101101111";
	Exp_in <= "01101001110000001101110111110000000011100000110110000010000001100011110011000110010111000010100000100010101111100001011100011001";
	M_in <= "10000110110000000010001111101011101000100000111010100010001110100110011100010010100101101111101001101010100010010111100110001101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01011100010000001011001101001011000001010110001001100000101000110010001001010010000101000101110101000010100001011011110011111000") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=163234658096966421351996810315840651486, exp=65537, mod=257052728932580766975123005399696262839";
	REPORT "Expected output is 209214796095670048995874763830207185992, 10011101011001010100110111010110111100000100010100100010010010000000110111101001001000011011111101101111100010000000010001001000";
	N_in <= "01111010110011011101101000000010011001011010010010111001001000101000100010010011000010100101111000010101010111001000000011011110";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "11000001011000101000111000000110111101101110111110001001110111111000010001010011101101000110100001101110111101011100011010110111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "10011101011001010100110111010110111100000100010100100010010010000000110111101001001000011011111101101111100010000000010001001000") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=209214796095670048995874763830207185992, exp=116306583625094488219330164562281959393, mod=257052728932580766975123005399696262839";
	REPORT "Expected output is 163234658096966421351996810315840651486, 01111010110011011101101000000010011001011010010010111001001000101000100010010011000010100101111000010101010111001000000011011110";
	N_in <= "10011101011001010100110111010110111100000100010100100010010010000000110111101001001000011011111101101111100010000000010001001000";
	Exp_in <= "01010111011111111101010101001101011101110110101110011000110010100101011111101001100100010110101101100101110010010000111111100001";
	M_in <= "11000001011000101000111000000110111101101110111110001001110111111000010001010011101101000110100001101110111101011100011010110111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01111010110011011101101000000010011001011010010010111001001000101000100010010011000010100101111000010101010111001000000011011110") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=143255536011528045391679156626753187552, exp=65537, mod=207856675875925324898784024365617151797";
	REPORT "Expected output is 97871591650611460179669960477144957034, 01001001101000010110001000000110001010001010010010010011100110100011101100111110001001100101011101000011001100101100000001101010";
	N_in <= "01101011110001100000001100111101000011100011110000010101011010010001110100111101010010011001110101100000010101011110111011100000";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10011100010111111011110101010111110011011010110000001010010111010000101101000000010110010111001100010100001001000111111100110101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01001001101000010110001000000110001010001010010010010011100110100011101100111110001001100101011101000011001100101100000001101010") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=97871591650611460179669960477144957034, exp=29638534508148407148928294312944902273, mod=207856675875925324898784024365617151797";
	REPORT "Expected output is 143255536011528045391679156626753187552, 01101011110001100000001100111101000011100011110000010101011010010001110100111101010010011001110101100000010101011110111011100000";
	N_in <= "01001001101000010110001000000110001010001010010010010011100110100011101100111110001001100101011101000011001100101100000001101010";
	Exp_in <= "00010110010011000010110010010010100101011001100000111111100011001000010100010101111111001100111100001100010010001010000010000001";
	M_in <= "10011100010111111011110101010111110011011010110000001010010111010000101101000000010110010111001100010100001001000111111100110101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01101011110001100000001100111101000011100011110000010101011010010001110100111101010010011001110101100000010101011110111011100000") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=129712307644364713188360756130267298158, exp=65537, mod=182542455999888314602731941240641923331";
	REPORT "Expected output is 146328742171449242480453944233531823163, 01101110000101011110010000000000001001011100010101101111111101111001101000001011100110000010001000111011010000000101010000111011";
	N_in <= "01100001100101011010111010000110110100111000010001100000101100010100100001100100011101111011010101001000001100000111100101101110";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10001001010101000110010111110001010011010010100110110111110011111001110011100101000111011011000001101110010100111010100100000011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01101110000101011110010000000000001001011100010101101111111101111001101000001011100110000010001000111011010000000101010000111011") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=146328742171449242480453944233531823163, exp=66778390567119678018268720068219394673, mod=182542455999888314602731941240641923331";
	REPORT "Expected output is 129712307644364713188360756130267298158, 01100001100101011010111010000110110100111000010001100000101100010100100001100100011101111011010101001000001100000111100101101110";
	N_in <= "01101110000101011110010000000000001001011100010101101111111101111001101000001011100110000010001000111011010000000101010000111011";
	Exp_in <= "00110010001111010000110011011010000111001001011101100001011000100110000011010111001011001110010100000010000001000101101001110001";
	M_in <= "10001001010101000110010111110001010011010010100110110111110011111001110011100101000111011011000001101110010100111010100100000011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01100001100101011010111010000110110100111000010001100000101100010100100001100100011101111011010101001000001100000111100101101110") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=90824878922666057384510049407850274714, exp=65537, mod=207405244049607743820860963498302134473";
	REPORT "Expected output is 88440021935079339884916747343563624727, 01000010100010001110110110111100001011101111111000100001111000000111000000000001001110001110110100101100000101001001000100010111";
	N_in <= "01000100010101000011110001000011010000011010000101111011010011000001101011110111101110001000110101111110011100000101111110011010";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10011100000010001100110000001001000110001101000010111011010101010000110111010001001011011001101011101110100100000101100011001001";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01000010100010001110110110111100001011101111111000100001111000000111000000000001001110001110110100101100000101001001000100010111") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=88440021935079339884916747343563624727, exp=43910276045414154482732384667249358973, mod=207405244049607743820860963498302134473";
	REPORT "Expected output is 90824878922666057384510049407850274714, 01000100010101000011110001000011010000011010000101111011010011000001101011110111101110001000110101111110011100000101111110011010";
	N_in <= "01000010100010001110110110111100001011101111111000100001111000000111000000000001001110001110110100101100000101001001000100010111";
	Exp_in <= "00100001000010001100111111000001110000010100101000110111110011000110100111000000010001000000101010110110110111110011100001111101";
	M_in <= "10011100000010001100110000001001000110001101000010111011010101010000110111010001001011011001101011101110100100000101100011001001";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01000100010101000011110001000011010000011010000101111011010011000001101011110111101110001000110101111110011100000101111110011010") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=161089105713639695570858797630103598343, exp=65537, mod=198637559406150265061528981782036962431";
	REPORT "Expected output is 8685567045391745169113773817473234444, 00000110100010001100011110000100100000100011000110001000110101001100100000010001100100111101100011110110110111110111011000001100";
	N_in <= "01111001001100001010001000011100000100100111001111101001111010001110000101101100100100110111110001011100010011011011010100000111";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10010101011100000011001111001110110010001101000111001100111010011000001001101111010000010101101100100111011010110101110001111111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "00000110100010001100011110000100100000100011000110001000110101001100100000010001100100111101100011110110110111110111011000001100") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=8685567045391745169113773817473234444, exp=181618930294876728690227506593114580673, mod=198637559406150265061528981782036962431";
	REPORT "Expected output is 161089105713639695570858797630103598343, 01111001001100001010001000011100000100100111001111101001111010001110000101101100100100110111110001011100010011011011010100000111";
	N_in <= "00000110100010001100011110000100100000100011000110001000110101001100100000010001100100111101100011110110110111110111011000001100";
	Exp_in <= "10001000101000101000100010011100000111110111110111000100100000111100110101111000111010110111101010100001001011110110011011000001";
	M_in <= "10010101011100000011001111001110110010001101000111001100111010011000001001101111010000010101101100100111011010110101110001111111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01111001001100001010001000011100000100100111001111101001111010001110000101101100100100110111110001011100010011011011010100000111") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=93221943264439933807802501486049021221, exp=65537, mod=222822424945745224760747010232056943463";
	REPORT "Expected output is 91702338258661188521183401408947963164, 01000100111111010011101001011001000111010010000001001110101000000000001010001110101100011110001001000100101010100100010100011100";
	N_in <= "01000110001000011110010010101000110011001111111100000100010011011111101101001011101111011111010010101000000010001100110100100101";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10100111101000100000100110111101100010100011010010010001110000111001010110001000011010101010100011010011001101100001001101100111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01000100111111010011101001011001000111010010000001001110101000000000001010001110101100011110001001000100101010100100010100011100") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=91702338258661188521183401408947963164, exp=110161731398554877687758338167710446353, mod=222822424945745224760747010232056943463";
	REPORT "Expected output is 93221943264439933807802501486049021221, 01000110001000011110010010101000110011001111111100000100010011011111101101001011101111011111010010101000000010001100110100100101";
	N_in <= "01000100111111010011101001011001000111010010000001001110101000000000001010001110101100011110001001000100101010100100010100011100";
	Exp_in <= "01010010111000000110000010110010011011011010111010111001110011110001110000100011100100101000001101101011011111000111001100010001";
	M_in <= "10100111101000100000100110111101100010100011010010010001110000111001010110001000011010101010100011010011001101100001001101100111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01000110001000011110010010101000110011001111111100000100010011011111101101001011101111011111010010101000000010001100110100100101") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=127634532801663317500488586413924027466, exp=65537, mod=172524665518916293003281099321502960339";
	REPORT "Expected output is 1760822805980569757756709938677643042, 00000001010100110001111101000100010111001101000001011001010001000000110001010001011011011101001100111101001101110111011100100010";
	N_in <= "01100000000001011000010001010001010101011000011101011101110100101011100010111100100110000010011110110110011101100000110001001010";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10000001110010110000101010111101000001101111101101100100001101100100010110001000101011000010010001111100000101011000101011010011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "00000001010100110001111101000100010111001101000001011001010001000000110001010001011011011101001100111101001101110111011100100010") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=1760822805980569757756709938677643042, exp=19325015938696682876130765886932492281, mod=172524665518916293003281099321502960339";
	REPORT "Expected output is 127634532801663317500488586413924027466, 01100000000001011000010001010001010101011000011101011101110100101011100010111100100110000010011110110110011101100000110001001010";
	N_in <= "00000001010100110001111101000100010111001101000001011001010001000000110001010001011011011101001100111101001101110111011100100010";
	Exp_in <= "00001110100010011101110011011001000100011010100000100101001011110111001100101101000010101001100100000111110010011001111111111001";
	M_in <= "10000001110010110000101010111101000001101111101101100100001101100100010110001000101011000010010001111100000101011000101011010011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01100000000001011000010001010001010101011000011101011101110100101011100010111100100110000010011110110110011101100000110001001010") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=134912623839323569481388422500950988202, exp=65537, mod=193317154930841576962082455216025435137";
	REPORT "Expected output is 145528813779176429820634048369696139419, 01101101011110111101010001111100011000001001011010100111010100010110101100101001100011011111111000101100100101110110100010011011";
	N_in <= "01100101011111110011100111101001000101010000001111011111111000100000000100010111111000110000111001110111011101111101010110101010";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10010001011011111000011110011101010101011111111000010111000010101111000011110011010110000010101000101011110110101111110000000001";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01101101011110111101010001111100011000001001011010100111010100010110101100101001100011011111111000101100100101110110100010011011") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=145528813779176429820634048369696139419, exp=19061224272748192151386989406312603649, mod=193317154930841576962082455216025435137";
	REPORT "Expected output is 134912623839323569481388422500950988202, 01100101011111110011100111101001000101010000001111011111111000100000000100010111111000110000111001110111011101111101010110101010";
	N_in <= "01101101011110111101010001111100011000001001011010100111010100010110101100101001100011011111111000101100100101110110100010011011";
	Exp_in <= "00001110010101110000111011101010001001101001011001111101001100100001010011110011101010001100001000101111000101100010000000000001";
	M_in <= "10010001011011111000011110011101010101011111111000010111000010101111000011110011010110000010101000101011110110101111110000000001";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01100101011111110011100111101001000101010000001111011111111000100000000100010111111000110000111001110111011101111101010110101010") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=133918481981842647051456135726411562113, exp=65537, mod=244525080833792013422574231312568015021";
	REPORT "Expected output is 243182735601533630516857329277366536577, 10110110111100110100101010001111000011010100110110001111001110010100110100101011010000100001010101011001010010011000100110000001";
	N_in <= "01100100101111111100001011101110110000001001100000110011010011001010100001010001101001110010110110010111011011000011110010000001";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10110111111101011101000101001001110110100100001010101111010100011111111000000100000000001101011101011001011111011101100010101101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "10110110111100110100101010001111000011010100110110001111001110010100110100101011010000100001010101011001010010011000100110000001") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=243182735601533630516857329277366536577, exp=77095713036432005868973642271493773121, mod=244525080833792013422574231312568015021";
	REPORT "Expected output is 133918481981842647051456135726411562113, 01100100101111111100001011101110110000001001100000110011010011001010100001010001101001110010110110010111011011000011110010000001";
	N_in <= "10110110111100110100101010001111000011010100110110001111001110010100110100101011010000100001010101011001010010011000100110000001";
	Exp_in <= "00111010000000000001100000011111100101111110000001000100100100001100011111010101000011000000000000111010111000001101011101000001";
	M_in <= "10110111111101011101000101001001110110100100001010101111010100011111111000000100000000001101011101011001011111011101100010101101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01100100101111111100001011101110110000001001100000110011010011001010100001010001101001110010110110010111011011000011110010000001") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=100920415182223406911780227792056066017, exp=65537, mod=221350269456308153845719435431166841213";
	REPORT "Expected output is 196780487042451605393567648295175643542, 10010100000010101000101100010010001101011101001000111110011111111110010001111000101010111000000101111010111100001110000110010110";
	N_in <= "01001011111011001001000010100001001101110000000101101110100010101100101010101110010110010110010010110010111111111001111111100001";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10100110100001101000001011011110111100101000111010110101111101111000011111110011100111101111110001001000001110111001000101111101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "10010100000010101000101100010010001101011101001000111110011111111110010001111000101010111000000101111010111100001110000110010110") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=196780487042451605393567648295175643542, exp=97055424311403803964611750436841766657, mod=221350269456308153845719435431166841213";
	REPORT "Expected output is 100920415182223406911780227792056066017, 01001011111011001001000010100001001101110000000101101110100010101100101010101110010110010110010010110010111111111001111111100001";
	N_in <= "10010100000010101000101100010010001101011101001000111110011111111110010001111000101010111000000101111010111100001110000110010110";
	Exp_in <= "01001001000001000011000111011110000011111111110100000011010001011100000111111101101101000011010111100110100101001011111100000001";
	M_in <= "10100110100001101000001011011110111100101000111010110101111101111000011111110011100111101111110001001000001110111001000101111101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01001011111011001001000010100001001101110000000101101110100010101100101010101110010110010110010010110010111111111001111111100001") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=162105959002765637930733811173896691455, exp=65537, mod=175915649338747166208470885449927869613";
	REPORT "Expected output is 139155790507188352042418866495276201848, 01101000101100000110111000101101110111000010010011011010110011100101001111000001001010110010100001111001101010000011011101111000";
	N_in <= "01111001111101000111100011011000111110000110001110101011111100100101000100100111110001011011010010101010101110110001111011111111";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10000100010110000001111100100110000101000001100001111111101100000101110111010110100111010111001000011100110110011100010010101101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01101000101100000110111000101101110111000010010011011010110011100101001111000001001010110010100001111001101010000011011101111000") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=139155790507188352042418866495276201848, exp=116299149166118352370661293355492836481, mod=175915649338747166208470885449927869613";
	REPORT "Expected output is 162105959002765637930733811173896691455, 01111001111101000111100011011000111110000110001110101011111100100101000100100111110001011011010010101010101110110001111011111111";
	N_in <= "01101000101100000110111000101101110111000010010011011010110011100101001111000001001010110010100001111001101010000011011101111000";
	Exp_in <= "01010111011111100110011011000001011001101110000110110111011010000000100111110001111000001101001110001011000000100000010010000001";
	M_in <= "10000100010110000001111100100110000101000001100001111111101100000101110111010110100111010111001000011100110110011100010010101101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01111001111101000111100011011000111110000110001110101011111100100101000100100111110001011011010010101010101110110001111011111111") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=169640536599918224955249115817138250639, exp=65537, mod=199194597955002668190107968515588196087";
	REPORT "Expected output is 88715816422201329258064073060667462625, 01000010101111100000101101110100000000001111101001110010100101100001111101011100101011101000100110011100001010011001001111100001";
	N_in <= "01111111100111111001010000110100001110101111000010101011000000010100011011000111010011101000000001111000100000001110001110001111";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10010101110110110111101111101101101110100000100100101110010011101011111111110011000100011100111000011010010001111000011011110111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01000010101111100000101101110100000000001111101001110010100101100001111101011100101011101000100110011100001010011001001111100001") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=88715816422201329258064073060667462625, exp=65621120433472810801879544338430360993, mod=199194597955002668190107968515588196087";
	REPORT "Expected output is 169640536599918224955249115817138250639, 01111111100111111001010000110100001110101111000010101011000000010100011011000111010011101000000001111000100000001110001110001111";
	N_in <= "01000010101111100000101101110100000000001111101001110010100101100001111101011100101011101000100110011100001010011001001111100001";
	Exp_in <= "00110001010111100010101100000111011101111110000000001010011000110111011101101111101111100110000011010110011111001111110110100001";
	M_in <= "10010101110110110111101111101101101110100000100100101110010011101011111111110011000100011100111000011010010001111000011011110111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01111111100111111001010000110100001110101111000010101011000000010100011011000111010011101000000001111000100000001110001110001111") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=145572578565823642614397331624412698668, exp=65537, mod=188451372387738631582433584346609765251";
	REPORT "Expected output is 159311774607762645508944040991940385860, 01110111110110100101010011101011101010111100111011111100010000000010010101111010000010100110000010101111100100111001110001000100";
	N_in <= "01101101100001000100001001000001101001010000100110111111011001001100000100011101000110111100011011000001001111011101100000101100";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10001101110001100110101000000011011001000001010001011101111010101111001101110001101000011011000010100011100100000100101110000011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01110111110110100101010011101011101010111100111011111100010000000010010101111010000010100110000010101111100100111001110001000100") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=159311774607762645508944040991940385860, exp=78998497850196734937919420243434279873, mod=188451372387738631582433584346609765251";
	REPORT "Expected output is 145572578565823642614397331624412698668, 01101101100001000100001001000001101001010000100110111111011001001100000100011101000110111100011011000001001111011101100000101100";
	N_in <= "01110111110110100101010011101011101010111100111011111100010000000010010101111010000010100110000010101111100100111001110001000100";
	Exp_in <= "00111011011011101000111010101000011001110011111011000110011011011010100011110011010110001000011011100000111110000001001111000001";
	M_in <= "10001101110001100110101000000011011001000001010001011101111010101111001101110001101000011011000010100011100100000100101110000011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01101101100001000100001001000001101001010000100110111111011001001100000100011101000110111100011011000001001111011101100000101100") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=148841961347667921326895815275312675983, exp=65537, mod=191898019277396571566977731419343411979";
	REPORT "Expected output is 66574649041872453527868538446945064230, 00110010000101011100111110011110100001101110111011100100101000100011010111001101001000101010101111111011111010100001010100100110";
	N_in <= "01101111111110011110101101000101110100010100011000000101000011011110011001110100010100000000100101101111010110010111110010001111";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10010000010111100011011011010011001010000001010110011011111101111011110000010110100100101111101000101001101010111101101100001011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "00110010000101011100111110011110100001101110111011100100101000100011010111001101001000101010101111111011111010100001010100100110") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=66574649041872453527868538446945064230, exp=77755342812628987466065822308881901873, mod=191898019277396571566977731419343411979";
	REPORT "Expected output is 148841961347667921326895815275312675983, 01101111111110011110101101000101110100010100011000000101000011011110011001110100010100000000100101101111010110010111110010001111";
	N_in <= "00110010000101011100111110011110100001101110111011100100101000100011010111001101001000101010101111111011111010100001010100100110";
	Exp_in <= "00111010011111110010001001100001110111101111110100011010100001110011010101100001000010110101000011100110000110111010100100110001";
	M_in <= "10010000010111100011011011010011001010000001010110011011111101111011110000010110100100101111101000101001101010111101101100001011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01101111111110011110101101000101110100010100011000000101000011011110011001110100010100000000100101101111010110010111110010001111") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=152924351631398877129203069757210809932, exp=65537, mod=284899033951435211130266243283506191373";
	REPORT "Expected output is 26491333971711071757281509514846017493, 00010011111011100000101110011011001010001011001011001011101111010001011000100110010111110000100110100001010111100001011111010101";
	N_in <= "01110011000011000010100010100111010101010001111100011110110001100101010010000001101111111001011100110000101100001101011001001100";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "11010110010101011000111011011101000111001100001000000001101011001010000011110101010100110100011100111010111000000101110000001101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "00010011111011100000101110011011001010001011001011001011101111010001011000100110010111110000100110100001010111100001011111010101") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=26491333971711071757281509514846017493, exp=180171893146637529180011746053852463937, mod=284899033951435211130266243283506191373";
	REPORT "Expected output is 152924351631398877129203069757210809932, 01110011000011000010100010100111010101010001111100011110110001100101010010000001101111111001011100110000101100001101011001001100";
	N_in <= "00010011111011100000101110011011001010001011001011001011101111010001011000100110010111110000100110100001010111100001011111010101";
	Exp_in <= "10000111100010111101100000101011100100011001001001000111101111111111111010011100111001100100000100101111010100111000001101000001";
	M_in <= "11010110010101011000111011011101000111001100001000000001101011001010000011110101010100110100011100111010111000000101110000001101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01110011000011000010100010100111010101010001111100011110110001100101010010000001101111111001011100110000101100001101011001001100") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=153699250002834601584677136791144568687, exp=65537, mod=233659187837269399573973084644251445987";
	REPORT "Expected output is 96164207072791911173816857966496046573, 01001000010110001000110101110111000011111001010000110101101000000100010001001000100001101011100011101101111001011101110111101101";
	N_in <= "01110011101000010110011000010111110100110000110110101010100101001011111000101110000001011111000101000000010001010001011101101111";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10101111110010010001111101100110111000110110001101110100101010010111000011001011011001100001011100101000001100101010101011100011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01001000010110001000110101110111000011111001010000110101101000000100010001001000100001101011100011101101111001011101110111101101") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=96164207072791911173816857966496046573, exp=125826633156124199179966596396815936033, mod=233659187837269399573973084644251445987";
	REPORT "Expected output is 153699250002834601584677136791144568687, 01110011101000010110011000010111110100110000110110101010100101001011111000101110000001011111000101000000010001010001011101101111";
	N_in <= "01001000010110001000110101110111000011111001010000110101101000000100010001001000100001101011100011101101111001011101110111101101";
	Exp_in <= "01011110101010010101001111111011101110000001111111101010110000000100111101110101111110000011111011101110101011101110101000100001";
	M_in <= "10101111110010010001111101100110111000110110001101110100101010010111000011001011011001100001011100101000001100101010101011100011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01110011101000010110011000010111110100110000110110101010100101001011111000101110000001011111000101000000010001010001011101101111") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=90433705321087480663210780013630059624, exp=65537, mod=197326791385053462287776461148218857119";
	REPORT "Expected output is 90170902292406843823174639973870785994, 01000011110101100100100010111001101101100011010001001100111010110001101110111100111101100011110000110111100000101101010111001010";
	N_in <= "01000100000010001110010111101010010001011111100100100011111110101011010101101000011000000101101100001101001001111111010001101000";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10010100011100111100000111110100011011000000010000000110111101111011100011000010101101110111000001010100010101100001011010011111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01000011110101100100100010111001101101100011010001001100111010110001101110111100111101100011110000110111100000101101010111001010") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=90170902292406843823174639973870785994, exp=117802321023852429977091988975366873473, mod=197326791385053462287776461148218857119";
	REPORT "Expected output is 90433705321087480663210780013630059624, 01000100000010001110010111101010010001011111100100100011111110101011010101101000011000000101101100001101001001111111010001101000";
	N_in <= "01000011110101100100100010111001101101100011010001001100111010110001101110111100111101100011110000110111100000101101010111001010";
	Exp_in <= "01011000100111111110011011011001100110011010011010101001110011110001101011000011000011100110011100101010110000101010000110000001";
	M_in <= "10010100011100111100000111110100011011000000010000000110111101111011100011000010101101110111000001010100010101100001011010011111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01000100000010001110010111101010010001011111100100100011111110101011010101101000011000000101101100001101001001111111010001101000") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=166857464301849188265314074580067827379, exp=65537, mod=183996335498353573095333378608267500559";
	REPORT "Expected output is 36742512848218808970092659623138262743, 00011011101001000101100110111111001000001110111100011111101111000000110011111001010011001000011000110110000101010111111011010111";
	N_in <= "01111101100001111001010000100101010100000000100010001111010011101111100101010011000101111001000000011110111100000011111010110011";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10001010011011000110011110111100011101010001000001111111110010101111100110001000011011011010101001101100101110111001110000001111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "00011011101001000101100110111111001000001110111100011111101111000000110011111001010011001000011000110110000101010111111011010111") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=36742512848218808970092659623138262743, exp=102623221256257047948682500544973529977, mod=183996335498353573095333378608267500559";
	REPORT "Expected output is 166857464301849188265314074580067827379, 01111101100001111001010000100101010100000000100010001111010011101111100101010011000101111001000000011110111100000011111010110011";
	N_in <= "00011011101001000101100110111111001000001110111100011111101111000000110011111001010011001000011000110110000101010111111011010111";
	Exp_in <= "01001101001101001000001101110011011110000111001110011000010111100110101001011111011110111010001011001100110110000110001101111001";
	M_in <= "10001010011011000110011110111100011101010001000001111111110010101111100110001000011011011010101001101100101110111001110000001111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01111101100001111001010000100101010100000000100010001111010011101111100101010011000101111001000000011110111100000011111010110011") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=86527273016340747463799613805957292284, exp=65537, mod=267436384001867615236177062946100009071";
	REPORT "Expected output is 4152667937977029627279567889007957076, 00000011000111111100011001010110001101111101100100101000010111110011111000011111010001000100011000010101111110001101010001010100";
	N_in <= "01000001000110001000101111101110101100000000011111001101010101100011011111010101000010101111111000001100010100010010000011111100";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "11001001001100100101111110111111100100000101111110010101101100010010101011100001010011001110010100000010101111001101100001101111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "00000011000111111100011001010110001101111101100100101000010111110011111000011111010001000100011000010101111110001101010001010100") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=4152667937977029627279567889007957076, exp=257495815598850242980319948614747365185, mod=267436384001867615236177062946100009071";
	REPORT "Expected output is 86527273016340747463799613805957292284, 01000001000110001000101111101110101100000000011111001101010101100011011111010101000010101111111000001100010100010010000011111100";
	N_in <= "00000011000111111100011001010110001101111101100100101000010111110011111000011111010001000100011000010101111110001101010001010100";
	Exp_in <= "11000001101101111110001111100010111100010110001001100111000101011010111000001101011110111100100101101000011101010001111101000001";
	M_in <= "11001001001100100101111110111111100100000101111110010101101100010010101011100001010011001110010100000010101111001101100001101111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01000001000110001000101111101110101100000000011111001101010101100011011111010101000010101111111000001100010100010010000011111100") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=121662052396835691967005993570708793081, exp=65537, mod=196731377532880914557844424081696334363";
	REPORT "Expected output is 113912343486356712974870877920718940577, 01010101101100101011100000100110011000000011101101110000000111010011111101000001001001010101010011110010101001101110100110100001";
	N_in <= "01011011100001110100001001001100100011101001100100011000101101000101011111010100001100000010000000100100101001001010011011111001";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10010100000000010001010111001001000011100011000101100001100111100001010000010101111110111100010001010001000111111010001000011011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01010101101100101011100000100110011000000011101101110000000111010011111101000001001001010101010011110010101001101110100110100001") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=113912343486356712974870877920718940577, exp=113910700569758030693755000099675214441, mod=196731377532880914557844424081696334363";
	REPORT "Expected output is 121662052396835691967005993570708793081, 01011011100001110100001001001100100011101001100100011000101101000101011111010100001100000010000000100100101001001010011011111001";
	N_in <= "01010101101100101011100000100110011000000011101101110000000111010011111101000001001001010101010011110010101001101110100110100001";
	Exp_in <= "01010101101100100110011100100101110110100110010011110111011001100000000110011000011011010011100011000000111110101001001001101001";
	M_in <= "10010100000000010001010111001001000011100011000101100001100111100001010000010101111110111100010001010001000111111010001000011011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01011011100001110100001001001100100011101001100100011000101101000101011111010100001100000010000000100100101001001010011011111001") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=86989139211378037676316071605009903497, exp=65537, mod=195347412942832780479598643425274334827";
	REPORT "Expected output is 119895152452813224471817881321061560241, 01011010001100101111011101100111111011011011100010101110011110001011100110110110100110100001010000011100010010010010111110110001";
	N_in <= "01000001011100010111111110110001101001001001100001001000101100011111100000000001000101011011100000011111011000111110111110001001";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10010010111101101000101100010000000110110100110110101010011110110011100001110011011110010011010001111010001101011000111001101011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01011010001100101111011101100111111011011011100010101110011110001011100110110110100110100001010000011100010010010010111110110001") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=119895152452813224471817881321061560241, exp=9046483639493682773137370833494395873, mod=195347412942832780479598643425274334827";
	REPORT "Expected output is 86989139211378037676316071605009903497, 01000001011100010111111110110001101001001001100001001000101100011111100000000001000101011011100000011111011000111110111110001001";
	N_in <= "01011010001100101111011101100111111011011011100010101110011110001011100110110110100110100001010000011100010010010010111110110001";
	Exp_in <= "00000110110011100100101000010100010111011101111101010011111001000001101001101101001110011010000000000001001000101100101111100001";
	M_in <= "10010010111101101000101100010000000110110100110110101010011110110011100001110011011110010011010001111010001101011000111001101011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01000001011100010111111110110001101001001001100001001000101100011111100000000001000101011011100000011111011000111110111110001001") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=148875969347815660350369849701071046314, exp=65537, mod=190168773485728868850383357234743879031";
	REPORT "Expected output is 62660687505308883530459386830636174237, 00101111001001000000001001101010101011001110001100111111111101011101000111110001111011001010100000000001011101111100101110011101";
	N_in <= "01110000000000000111011111111111001000000011111111101110000100100010011001111110101010110100010100001010110101111100011010101010";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10001111000100010010110001101100101111110101111100101100011100110110001101110001101100001011000011110111100001000010010101110111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "00101111001001000000001001101010101011001110001100111111111101011101000111110001111011001010100000000001011101111100101110011101") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=62660687505308883530459386830636174237, exp=67621238343400301440197569386348068161, mod=190168773485728868850383357234743879031";
	REPORT "Expected output is 148875969347815660350369849701071046314, 01110000000000000111011111111111001000000011111111101110000100100010011001111110101010110100010100001010110101111100011010101010";
	N_in <= "00101111001001000000001001101010101011001110001100111111111101011101000111110001111011001010100000000001011101111100101110011101";
	Exp_in <= "00110010110111110110000001110100101010101111100000100100110010101100100100011110111010111101110111000001110001001011110101000001";
	M_in <= "10001111000100010010110001101100101111110101111100101100011100110110001101110001101100001011000011110111100001000010010101110111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01110000000000000111011111111111001000000011111111101110000100100010011001111110101010110100010100001010110101111100011010101010") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=85584314150133822438826175682412715156, exp=65537, mod=182039830930609931786609312357468796457";
	REPORT "Expected output is 129571219152728082471381848214417833955, 01100001011110101000001001010011101100111101110000110100111011111111011010100010000011001000011000101010101110011111111111100011";
	N_in <= "01000000011000101111000001111000100001111111011001110011000010110000001010111110101001101011100000111000000111101001110010010100";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10001000111100111001100010011101000001101111011110000100011100001000011110010011010100000111110101000010000101101111011000101001";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01100001011110101000001001010011101100111101110000110100111011111111011010100010000011001000011000101010101110011111111111100011") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=129571219152728082471381848214417833955, exp=157924143423712218387216877522766921613, mod=182039830930609931786609312357468796457";
	REPORT "Expected output is 85584314150133822438826175682412715156, 01000000011000101111000001111000100001111111011001110011000010110000001010111110101001101011100000111000000111101001110010010100";
	N_in <= "01100001011110101000001001010011101100111101110000110100111011111111011010100010000011001000011000101010101110011111111111100011";
	Exp_in <= "01110110110011110001010101101011110011001011101001111000010011110101111010111000100100010101011110111000101101011111111110001101";
	M_in <= "10001000111100111001100010011101000001101111011110000100011100001000011110010011010100000111110101000010000101101111011000101001";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01000000011000101111000001111000100001111111011001110011000010110000001010111110101001101011100000111000000111101001110010010100") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=121068503598395469756608908445314169830, exp=65537, mod=172372499163015502304899783616402524027";
	REPORT "Expected output is 132042697782175870710390559317494812274, 01100011010101100111111110100001100110101011011010001011101010100001011001100011010101111000000000011001000101110100111001110010";
	N_in <= "01011011000101001111001000010101011110100110011100110011001011110000100110000101110000100111010110001001000111111011101111100110";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10000001101011011011110001011011100110010101111101101001110100111010100101100010111101010101111011001001111000111000011101111011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01100011010101100111111110100001100110101011011010001011101010100001011001100011010101111000000000011001000101110100111001110010") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=132042697782175870710390559317494812274, exp=69985806952235828546567207443095995633, mod=172372499163015502304899783616402524027";
	REPORT "Expected output is 121068503598395469756608908445314169830, 01011011000101001111001000010101011110100110011100110011001011110000100110000101110000100111010110001001000111111011101111100110";
	N_in <= "01100011010101100111111110100001100110101011011010001011101010100001011001100011010101111000000000011001000101110100111001110010";
	Exp_in <= "00110100101001101100011010110000011001100100000001100000001000011111011100100100000100000100001000101011011110011100010011110001";
	M_in <= "10000001101011011011110001011011100110010101111101101001110100111010100101100010111101010101111011001001111000111000011101111011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01011011000101001111001000010101011110100110011100110011001011110000100110000101110000100111010110001001000111111011101111100110") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=133604485749493167591551218804947276766, exp=65537, mod=274456619968110053023589940368633048249";
	REPORT "Expected output is 21673033971893824475753251772539407225, 00010000010011100001001100010011001010101101000110110110010011010001011001011100101101110111011000000111001100010000101101111001";
	N_in <= "01100100100000110100100110111001000111100111001000000011111000011101010001000111011110101110110111100101101000011101001111011110";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "11001110011110100110110000011010110000000100011011001100111100000000010101110111111010101000000000001110001001010010110010111001";
	wait for 33409 * clk_period;
	ASSERT(C_out = "00010000010011100001001100010011001010101101000110110110010011010001011001011100101101110111011000000111001100010000101101111001") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=21673033971893824475753251772539407225, exp=33745387242367377283869717967108222793, mod=274456619968110053023589940368633048249";
	REPORT "Expected output is 133604485749493167591551218804947276766, 01100100100000110100100110111001000111100111001000000011111000011101010001000111011110101110110111100101101000011101001111011110";
	N_in <= "00010000010011100001001100010011001010101101000110110110010011010001011001011100101101110111011000000111001100010000101101111001";
	Exp_in <= "00011001011000110010000000001011101000011111110010010010100100000101010001000010110110010110011011011000011011101010111101001001";
	M_in <= "11001110011110100110110000011010110000000100011011001100111100000000010101110111111010101000000000001110001001010010110010111001";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01100100100000110100100110111001000111100111001000000011111000011101010001000111011110101110110111100101101000011101001111011110") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=114757702792810332475522532486323700909, exp=65537, mod=209337289174751424503619704190096518083";
	REPORT "Expected output is 129606521629176841147012569074047709103, 01100001100000010100111011011111100110010101100110111010110101011000110000000010010000110011000000001011110100001110111110101111";
	N_in <= "01010110010101011000011110010100111001100100011100100101010000111101001000110101010110101101011000010110111110010000010010101101";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10011101011111001110010100110110111101010110000100101100001011010011011111010001000011001001000101010010000000100010101111000011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01100001100000010100111011011111100110010101100110111010110101011000110000000010010000110011000000001011110100001110111110101111") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=129606521629176841147012569074047709103, exp=174651636441964972083117575822167320305, mod=209337289174751424503619704190096518083";
	REPORT "Expected output is 114757702792810332475522532486323700909, 01010110010101011000011110010100111001100100011100100101010000111101001000110101010110101101011000010110111110010000010010101101";
	N_in <= "01100001100000010100111011011111100110010101100110111010110101011000110000000010010000110011000000001011110100001110111110101111";
	Exp_in <= "10000011011001001010111010000000010110011101110101000110110010001111101110111101000001110010000111010011011000010010011011110001";
	M_in <= "10011101011111001110010100110110111101010110000100101100001011010011011111010001000011001001000101010010000000100010101111000011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01010110010101011000011110010100111001100100011100100101010000111101001000110101010110101101011000010110111110010000010010101101") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=165430981043216411480404357894779276685, exp=65537, mod=200239132257456490290299447435093786963";
	REPORT "Expected output is 43281167004392969703106996670939916316, 00100000100011111010011001001001010100000100111110101010101000010010101000011000010000001000010000000010110000011110100000011100";
	N_in <= "01111100011101001101100100010111010100010101000000001111011111001001011011010111101101000110000100111110110100011000110110001101";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10010110101001001010011101110010001000011111000110010101001110110000110101001110001000100010010101111011001100101100000101010011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "00100000100011111010011001001001010100000100111110101010101000010010101000011000010000001000010000000010110000011110100000011100") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=43281167004392969703106996670939916316, exp=134356403281953578803583500153494112769, mod=200239132257456490290299447435093786963";
	REPORT "Expected output is 165430981043216411480404357894779276685, 01111100011101001101100100010111010100010101000000001111011111001001011011010111101101000110000100111110110100011000110110001101";
	N_in <= "00100000100011111010011001001001010100000100111110101010101000010010101000011000010000001000010000000010110000011110100000011100";
	Exp_in <= "01100101000101000001101000011110101001001101001111111010101010111010001010010000011110000001010011000100010100110000101000000001";
	M_in <= "10010110101001001010011101110010001000011111000110010101001110110000110101001110001000100010010101111011001100101100000101010011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01111100011101001101100100010111010100010101000000001111011111001001011011010111101101000110000100111110110100011000110110001101") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=113251135016392116067999548819039551951, exp=65537, mod=170823664564573541048918956028446711073";
	REPORT "Expected output is 61295625658127882134418451795594181946, 00101110000111010001101110101011111000100101011101001101001110010100111100010101111010000001111011111000100110111111110100111010";
	N_in <= "01010101001100110110000000001110001011100111000011011111010110101001001001100010011010100001101101011110001011111000000111001111";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10000000100000110111000011101010100101011101010011011110100001011110110001101110111000011110011011101111101001010001110100100001";
	wait for 33409 * clk_period;
	ASSERT(C_out = "00101110000111010001101110101011111000100101011101001101001110010100111100010101111010000001111011111000100110111111110100111010") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=61295625658127882134418451795594181946, exp=36788458453459739620042196154592528649, mod=170823664564573541048918956028446711073";
	REPORT "Expected output is 113251135016392116067999548819039551951, 01010101001100110110000000001110001011100111000011011111010110101001001001100010011010100001101101011110001011111000000111001111";
	N_in <= "00101110000111010001101110101011111000100101011101001101001110010100111100010101111010000001111011111000100110111111110100111010";
	Exp_in <= "00011011101011010011001100001010001100100100111001101111110000111000000010111101100111100110110110010110011100000000100100001001";
	M_in <= "10000000100000110111000011101010100101011101010011011110100001011110110001101110111000011110011011101111101001010001110100100001";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01010101001100110110000000001110001011100111000011011111010110101001001001100010011010100001101101011110001011111000000111001111") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=167466789591625782731611274151982261933, exp=65537, mod=174762125637185202227882446992458465377";
	REPORT "Expected output is 138236350903369394510498782233868573067, 01100111111111110101101001001110100001111000000001100000010101111000111101101000000111111011001110010010011110110001100110001011";
	N_in <= "01111101111111001110111000110011101101010001001000000011101010010011101000011110010011110110010000110001100100111110011010101101";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10000011011110011111011000001010000011100101010000001001100110111100000111101100101001111001100000110111100001010100000001100001";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01100111111111110101101001001110100001111000000001100000010101111000111101101000000111111011001110010010011110110001100110001011") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=138236350903369394510498782233868573067, exp=100499488701256326816123394302589037057, mod=174762125637185202227882446992458465377";
	REPORT "Expected output is 167466789591625782731611274151982261933, 01111101111111001110111000110011101101010001001000000011101010010011101000011110010011110110010000110001100100111110011010101101";
	N_in <= "01100111111111110101101001001110100001111000000001100000010101111000111101101000000111111011001110010010011110110001100110001011";
	Exp_in <= "01001011100110110111111101011010000110010001001101001010110010100010001011100000001110101100011000111011101000000110101000000001";
	M_in <= "10000011011110011111011000001010000011100101010000001001100110111100000111101100101001111001100000110111100001010100000001100001";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01111101111111001110111000110011101101010001001000000011101010010011101000011110010011110110010000110001100100111110011010101101") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=87236941637304974756486416226129652421, exp=65537, mod=225843539335348999348043362436683134869";
	REPORT "Expected output is 168902057209521497338464825565224376801, 01111111000100010101101001011011111001110110011010000100001100010010100110110110110111001111011000010001011000000001100111100001";
	N_in <= "01000001101000010011100101001011111110101011111010100111011011111001001111010010101111011100110000010011100000011010101011000101";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10101001111001111110001000101110000011011110110111001001001101001000010101101100011011110011010010001101011001111111011110010101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01111111000100010101101001011011111001110110011010000100001100010010100110110110110111001111011000010001011000000001100111100001") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=168902057209521497338464825565224376801, exp=107930171536431796591178952649834657313, mod=225843539335348999348043362436683134869";
	REPORT "Expected output is 87236941637304974756486416226129652421, 01000001101000010011100101001011111110101011111010100111011011111001001111010010101111011100110000010011100000011010101011000101";
	N_in <= "01111111000100010101101001011011111001110110011010000100001100010010100110110110110111001111011000010001011000000001100111100001";
	Exp_in <= "01010001001100101001100001001101000110100010101100000001011011111110100000110100100001011001000011011101010111100111011000100001";
	M_in <= "10101001111001111110001000101110000011011110110111001001001101001000010101101100011011110011010010001101011001111111011110010101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01000001101000010011100101001011111110101011111010100111011011111001001111010010101111011100110000010011100000011010101011000101") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=129221657295404037574021711945125721644, exp=65537, mod=227636589678176624737452402871879779479";
	REPORT "Expected output is 35081478336896887758341338200602986419, 00011010011001000111001001101100000111100000110000100011011000001001011000110001000101100011001001110001101011100100011110110011";
	N_in <= "01100001001101110010111110011000110001010111100110111010101100010001101000001001011010010110001001010011111100011111011000101100";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10101011010000010011011001100011000111101000010001011011011111101000110110100000111100000011000111000110101001101100010010010111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "00011010011001000111001001101100000111100000110000100011011000001001011000110001000101100011001001110001101011100100011110110011") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=35081478336896887758341338200602986419, exp=2219506245393516075703870490669060345, mod=227636589678176624737452402871879779479";
	REPORT "Expected output is 129221657295404037574021711945125721644, 01100001001101110010111110011000110001010111100110111010101100010001101000001001011010010110001001010011111100011111011000101100";
	N_in <= "00011010011001000111001001101100000111100000110000100011011000001001011000110001000101100011001001110001101011100100011110110011";
	Exp_in <= "00000001101010110111011000011011010010110100110111100001000100100101111100111110001000111011100011011010000000011001000011111001";
	M_in <= "10101011010000010011011001100011000111101000010001011011011111101000110110100000111100000011000111000110101001101100010010010111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01100001001101110010111110011000110001010111100110111010101100010001101000001001011010010110001001010011111100011111011000101100") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=93032806917345403385496193805259654666, exp=65537, mod=220915454521144462227553499198418902503";
	REPORT "Expected output is 83405139601179821116294329382504901871, 00111110101111110011111011011110110100000101111010110101111101011001110010101111111000000101010101011110100110100010110011101111";
	N_in <= "01000101111111010111011110000100011110110010100101010010001100101001000010101000111010000100110111000010100001000100011000001010";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10100110001100101100010011010110111001001100111011001101101010010010111100000011010011101000011000001011101001001101110111100111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "00111110101111110011111011011110110100000101111010110101111101011001110010101111111000000101010101011110100110100010110011101111") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=83405139601179821116294329382504901871, exp=51213337512241143338004566464445705353, mod=220915454521144462227553499198418902503";
	REPORT "Expected output is 93032806917345403385496193805259654666, 01000101111111010111011110000100011110110010100101010010001100101001000010101000111010000100110111000010100001000100011000001010";
	N_in <= "00111110101111110011111011011110110100000101111010110101111101011001110010101111111000000101010101011110100110100010110011101111";
	Exp_in <= "00100110100001110101010001111100101000001111010010010100010100111101110111110111100010100100110000001001100100100110110010001001";
	M_in <= "10100110001100101100010011010110111001001100111011001101101010010010111100000011010011101000011000001011101001001101110111100111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01000101111111010111011110000100011110110010100101010010001100101001000010101000111010000100110111000010100001000100011000001010") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=97647624986562465329317246022064063288, exp=65537, mod=170376124650059692302928940764746875363";
	REPORT "Expected output is 126286059366916285096059952336555117736, 01011111000000011100111101110001101111100110000111010100101111101111011011011011011001000101110100111101011100101000110010101000";
	N_in <= "01001001011101100011111110011101011011101110110100010010001000110011111111101010100110010111001000000101101011001100001100111000";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10000000001011010011111101111110101101100011111101011111110010101000111000001100111011111011000110010111100101100000000111100011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01011111000000011100111101110001101111100110000111010100101111101111011011011011011001000101110100111101011100101000110010101000") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=126286059366916285096059952336555117736, exp=46799685611950113338064751568646177473, mod=170376124650059692302928940764746875363";
	REPORT "Expected output is 97647624986562465329317246022064063288, 01001001011101100011111110011101011011101110110100010010001000110011111111101010100110010111001000000101101011001100001100111000";
	N_in <= "01011111000000011100111101110001101111100110000111010100101111101111011011011011011001000101110100111101011100101000110010101000";
	Exp_in <= "00100011001101010100101010100101101100011100011000000010101101011001001110011101110110001101010000011100011101100000001011000001";
	M_in <= "10000000001011010011111101111110101101100011111101011111110010101000111000001100111011111011000110010111100101100000000111100011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01001001011101100011111110011101011011101110110100010010001000110011111111101010100110010111001000000101101011001100001100111000") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=131147416515642893412630985167106455475, exp=65537, mod=171415913885036945633821271379370983853";
	REPORT "Expected output is 5553153113296698787854473536685552304, 00000100001011010111111110010110010001001100000110000100000110000100010111000000101011011000001011110000110010010011001010110000";
	N_in <= "01100010101010100001001011011011010110111101110010001100000001100001000010110111000110010001000000001010111110111011011110110011";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10000000111101011000000100001111111100100011100111100111000100100101101001011110011100001110100001111110011111100100000110101101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "00000100001011010111111110010110010001001100000110000100000110000100010111000000101011011000001011110000110010010011001010110000") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=5553153113296698787854473536685552304, exp=107033920197804017258875708329298954113, mod=171415913885036945633821271379370983853";
	REPORT "Expected output is 131147416515642893412630985167106455475, 01100010101010100001001011011011010110111101110010001100000001100001000010110111000110010001000000001010111110111011011110110011";
	N_in <= "00000100001011010111111110010110010001001100000110000100000110000100010111000000101011011000001011110000110010010011001010110000";
	Exp_in <= "01010000100001011111101110110010110100110101001101101000011101110110000110110001010100100100010010011110000111110000011110000001";
	M_in <= "10000000111101011000000100001111111100100011100111100111000100100101101001011110011100001110100001111110011111100100000110101101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01100010101010100001001011011011010110111101110010001100000001100001000010110111000110010001000000001010111110111011011110110011") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=93352691429873341459285693054896417079, exp=65537, mod=174770482091518834617139533444480828677";
	REPORT "Expected output is 31396861601783176929191607798479718353, 00010111100111101101000011001010101000001110010110100100010101110001000001001110010100010100111111100011011110000000011111010001";
	N_in <= "01000110001110110001001100001010101010001011010001101000010101011000101000010110111010110100011000011000010100011010100100110111";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10000011011110111001001000001011010101101000101010000000110000101111111001000010010100010000011000100011110101010000010100000101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "00010111100111101101000011001010101000001110010110100100010101110001000001001110010100010100111111100011011110000000011111010001") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=31396861601783176929191607798479718353, exp=9685618672755793006863876034299885569, mod=174770482091518834617139533444480828677";
	REPORT "Expected output is 93352691429873341459285693054896417079, 01000110001110110001001100001010101010001011010001101000010101011000101000010110111010110100011000011000010100011010100100110111";
	N_in <= "00010111100111101101000011001010101000001110010110100100010101110001000001001110010100010100111111100011011110000000011111010001";
	Exp_in <= "00000111010010010110000111011110100111101111110100101110000001001100010010000011001101100101010011110111011000101111100000000001";
	M_in <= "10000011011110111001001000001011010101101000101010000000110000101111111001000010010100010000011000100011110101010000010100000101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01000110001110110001001100001010101010001011010001101000010101011000101000010110111010110100011000011000010100011010100100110111") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=106387618117775449555072843817718323833, exp=65537, mod=210051512776609004203918952562644308967";
	REPORT "Expected output is 168739084726534070189168291788204591275, 01111110111100011111011100110001111110100000001110110000010000011100111100110101101100001101110110011001001000001100100010101011";
	N_in <= "01010000000010011000001010001011101110010001111100010100110111101100011100100100011111100000110101000010100110110001101001111001";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10011110000001100111001100101000001100010010010110001110000110101100100001111100000010101001001100011101101001010101001111100111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01111110111100011111011100110001111110100000001110110000010000011100111100110101101100001101110110011001001000001100100010101011") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=168739084726534070189168291788204591275, exp=46589083872023261382801122291202531521, mod=210051512776609004203918952562644308967";
	REPORT "Expected output is 106387618117775449555072843817718323833, 01010000000010011000001010001011101110010001111100010100110111101100011100100100011111100000110101000010100110110001101001111001";
	N_in <= "01111110111100011111011100110001111110100000001110110000010000011100111100110101101100001101110110011001001000001100100010101011";
	Exp_in <= "00100011000011001011101100101110000001101111100010010101011100010001100100110100010110011110111011101100000111100010000011000001";
	M_in <= "10011110000001100111001100101000001100010010010110001110000110101100100001111100000010101001001100011101101001010101001111100111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01010000000010011000001010001011101110010001111100010100110111101100011100100100011111100000110101000010100110110001101001111001") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=115528328906465421347117452505154314700, exp=65537, mod=178123323768742237134777495130072152701";
	REPORT "Expected output is 14486338350679677536132218645864001556, 00001010111001011111011110011111110000010010010110100001110111100010001011010101010101010100010001011000111010000011000000010100";
	N_in <= "01010110111010011111001001100001111010101100110110111000100110100100000000000000110100100111100111100010010111111110000111001100";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10000110000000010100110111100110110111011111000101111010010011101111101000001001111011101110000110110001000000111111101001111101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "00001010111001011111011110011111110000010010010110100001110111100010001011010101010101010100010001011000111010000011000000010100") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=14486338350679677536132218645864001556, exp=148082322538659872038062748942173518897, mod=178123323768742237134777495130072152701";
	REPORT "Expected output is 115528328906465421347117452505154314700, 01010110111010011111001001100001111010101100110110111000100110100100000000000000110100100111100111100010010111111110000111001100";
	N_in <= "00001010111001011111011110011111110000010010010110100001110111100010001011010101010101010100010001011000111010000011000000010100";
	Exp_in <= "01101111011001111001111000110000000101001100101110110000011010110010110101110011010111010100101101000101001000001011110000110001";
	M_in <= "10000110000000010100110111100110110111011111000101111010010011101111101000001001111011101110000110110001000000111111101001111101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01010110111010011111001001100001111010101100110110111000100110100100000000000000110100100111100111100010010111111110000111001100") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=128546278755025971076837868605050272066, exp=65537, mod=198370131366760057647013501598187185087";
	REPORT "Expected output is 56288968938165648761290790353681370995, 00101010010110001101110001101111110110010010101000110101100010000110010111111100110110100000011000101001100011011100111101110011";
	N_in <= "01100000101101010001110011011101001001001100101010100001011001110110111010010111010101100111001000101000000010010011100101000010";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10010101001111001011001010010110011000010111010100100111010010001101100011010101011110101111100011010011001101001110001110111111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "00101010010110001101110001101111110110010010101000110101100010000110010111111100110110100000011000101001100011011100111101110011") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=56288968938165648761290790353681370995, exp=175187549983144461979943965296563472497, mod=198370131366760057647013501598187185087";
	REPORT "Expected output is 128546278755025971076837868605050272066, 01100000101101010001110011011101001001001100101010100001011001110110111010010111010101100111001000101000000010010011100101000010";
	N_in <= "00101010010110001101110001101111110110010010101000110101100010000110010111111100110110100000011000101001100011011100111101110011";
	Exp_in <= "10000011110010111110010100010100001101011110000110010110110101000110100001000011011001001110110101000111100000100100100001110001";
	M_in <= "10010101001111001011001010010110011000010111010100100111010010001101100011010101011110101111100011010011001101001110001110111111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01100000101101010001110011011101001001001100101010100001011001110110111010010111010101100111001000101000000010010011100101000010") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=89267004892172012823271030719322226643, exp=65537, mod=199124812965268505113585587223215251741";
	REPORT "Expected output is 104509496073959389771722649366390902621, 01001110100111111100101111111010110101010110000111111000000010101000000100100000100000010100101111001111001100000000111101011101";
	N_in <= "01000011001010000011001100100100100100011101100011110110101101110101000011011010111000010101110111110010011001110111111111010011";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10010101110011100000101101000011010100101110110111011110011111110010010011101110001011001100000100111001100001001010000100011101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01001110100111111100101111111010110101010110000111111000000010101000000100100000100000010100101111001111001100000000111101011101") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=104509496073959389771722649366390902621, exp=172928097561961288410851111172910443713, mod=199124812965268505113585587223215251741";
	REPORT "Expected output is 89267004892172012823271030719322226643, 01000011001010000011001100100100100100011101100011110110101101110101000011011010111000010101110111110010011001110111111111010011";
	N_in <= "01001110100111111100101111111010110101010110000111111000000010101000000100100000100000010100101111001111001100000000111101011101";
	Exp_in <= "10000010000110001011110101111001010010110100010011011110110001000100100111010111001100011011001011001000110110010110110011000001";
	M_in <= "10010101110011100000101101000011010100101110110111011110011111110010010011101110001011001100000100111001100001001010000100011101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01000011001010000011001100100100100100011101100011110110101101110101000011011010111000010101110111110010011001110111111111010011") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=96902820348742501871409988685772628703, exp=65537, mod=172375998890493170635869297789266434643";
	REPORT "Expected output is 34764472254050610538055469097269604606, 00011010001001110110010011010000110101000110110001010001100110100110110110000101110101001001100110000010001011000011000011111110";
	N_in <= "01001000111001101100110111101001010000101010110011010001010010110011110111110000000011010010000111010011110001000010001011011111";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10000001101011100110100011101000010111101011111000101000111001001001111001100100001001011011101011110101100011100001101001010011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "00011010001001110110010011010000110101000110110001010001100110100110110110000101110101001001100110000010001011000011000011111110") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=34764472254050610538055469097269604606, exp=140826643462392012553903090415139844673, mod=172375998890493170635869297789266434643";
	REPORT "Expected output is 96902820348742501871409988685772628703, 01001000111001101100110111101001010000101010110011010001010010110011110111110000000011010010000111010011110001000010001011011111";
	N_in <= "00011010001001110110010011010000110101000110110001010001100110100110110110000101110101001001100110000010001011000011000011111110";
	Exp_in <= "01101001111100100011100110010111000011100100000001000001010011111011000001000100110000110111100110100000111111000111001001000001";
	M_in <= "10000001101011100110100011101000010111101011111000101000111001001001111001100100001001011011101011110101100011100001101001010011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01001000111001101100110111101001010000101010110011010001010010110011110111110000000011010010000111010011110001000010001011011111") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=89174818644703591002603786259083080590, exp=65537, mod=194897098142298662899482346320915367579";
	REPORT "Expected output is 13776246741884341492639181069824443201, 00001010010111010011010101100111100110110000100110001010100101001101000001010000111010111011100000100001010110100100001101000001";
	N_in <= "01000011000101100111001000000010100010110010111100010001110011111100000001111000011010110011110011010110000100001011001110001110";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10010010100111111101000011010100001111110110101000101000111110111001010001001101111001000011101101111100110011001000011010011011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "00001010010111010011010101100111100110110000100110001010100101001101000001010000111010111011100000100001010110100100001101000001") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=13776246741884341492639181069824443201, exp=57204946516704412376091771620055124001, mod=194897098142298662899482346320915367579";
	REPORT "Expected output is 89174818644703591002603786259083080590, 01000011000101100111001000000010100010110010111100010001110011111100000001111000011010110011110011010110000100001011001110001110";
	N_in <= "00001010010111010011010101100111100110110000100110001010100101001101000001010000111010111011100000100001010110100100001101000001";
	Exp_in <= "00101011000010010100010110011110010001101100111010111110000111000000111011011110001101101000010001100010001110010000100000100001";
	M_in <= "10010010100111111101000011010100001111110110101000101000111110111001010001001101111001000011101101111100110011001000011010011011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01000011000101100111001000000010100010110010111100010001110011111100000001111000011010110011110011010110000100001011001110001110") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=118331774880277334077242539021149112382, exp=65537, mod=287279728026516419963518043624318121647";
	REPORT "Expected output is 163644882903620607622399813668568275733, 01111011000111001101101110100111011001001110100101100001010111010000011001110011000000001101011000100001101100111001101100010101";
	N_in <= "01011001000001011101111011110000110001101000001011000111001110111101110011110101010000000010111001101010100101111000100000111110";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "11011000001000000001000000100100110101111010000100001011011001011100010110011111010110001011110010011110101011110011011010101111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01111011000111001101101110100111011001001110100101100001010111010000011001110011000000001101011000100001101100111001101100010101") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=163644882903620607622399813668568275733, exp=251642085338331447975463529012108373449, mod=287279728026516419963518043624318121647";
	REPORT "Expected output is 118331774880277334077242539021149112382, 01011001000001011101111011110000110001101000001011000111001110111101110011110101010000000010111001101010100101111000100000111110";
	N_in <= "01111011000111001101101110100111011001001110100101100001010111010000011001110011000000001101011000100001101100111001101100010101";
	Exp_in <= "10111101010100001000000010110011101101010000101001000101100001000100011011110111100101100001110100111000000010101010110111001001";
	M_in <= "11011000001000000001000000100100110101111010000100001011011001011100010110011111010110001011110010011110101011110011011010101111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01011001000001011101111011110000110001101000001011000111001110111101110011110101010000000010111001101010100101111000100000111110") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=120653453745836605323003298878166786541, exp=65537, mod=184897757648140267826328491935920982481";
	REPORT "Expected output is 45157183015557597314059792815223717735, 00100001111110001111010100000100010101011000101000011100010111010000010001101000000001100000100111001000010011111011111101100111";
	N_in <= "01011010110001010000001010001011110101101111011110000011101111110000001011011101000110100110000101101100100101011110000111101101";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10001011000110100000001101000111100010111101110111101100101001011011010101101111010010100000111010110101101011101000100111010001";
	wait for 33409 * clk_period;
	ASSERT(C_out = "00100001111110001111010100000100010101011000101000011100010111010000010001101000000001100000100111001000010011111011111101100111") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=45157183015557597314059792815223717735, exp=160919759841534165210009335531884082681, mod=184897757648140267826328491935920982481";
	REPORT "Expected output is 120653453745836605323003298878166786541, 01011010110001010000001010001011110101101111011110000011101111110000001011011101000110100110000101101100100101011110000111101101";
	N_in <= "00100001111110001111010100000100010101011000101000011100010111010000010001101000000001100000100111001000010011111011111101100111";
	Exp_in <= "01111001000100000000010010110110101010100010011001010101100111001100010011010111011001101011001101110000111001010111010111111001";
	M_in <= "10001011000110100000001101000111100010111101110111101100101001011011010101101111010010100000111010110101101011101000100111010001";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01011010110001010000001010001011110101101111011110000011101111110000001011011101000110100110000101101100100101011110000111101101") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=153660397790020801384664009444082169131, exp=65537, mod=178684616015241641884280350209520452791";
	REPORT "Expected output is 70907843034280174191676698452813170851, 00110101010110000101101010010011111001001000010111001111100111111011010111001000001100110101110100110000010110000100100010100011";
	N_in <= "01110011100110011110101010000111111101001100001101001110011101100011110111101011010001111100110010101110101001011011010100101011";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10000110011011010110011110111111000001011000101000011110110100100000000101001101110001001010000001011000000111000100010010110111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "00110101010110000101101010010011111001001000010111001111100111111011010111001000001100110101110100110000010110000100100010100011") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=70907843034280174191676698452813170851, exp=67842734643136819950205663987155519473, mod=178684616015241641884280350209520452791";
	REPORT "Expected output is 153660397790020801384664009444082169131, 01110011100110011110101010000111111101001100001101001110011101100011110111101011010001111100110010101110101001011011010100101011";
	N_in <= "00110101010110000101101010010011111001001000010111001111100111111011010111001000001100110101110100110000010110000100100010100011";
	Exp_in <= "00110011000010100000100100010001000000110001011001101101000101100110000110001000110001011111010010101000011101101100011111110001";
	M_in <= "10000110011011010110011110111111000001011000101000011110110100100000000101001101110001001010000001011000000111000100010010110111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01110011100110011110101010000111111101001100001101001110011101100011110111101011010001111100110010101110101001011011010100101011") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=113983681069878420564395489959401671234, exp=65537, mod=228444100611487427329574816502404255489";
	REPORT "Expected output is 191823984475670677583965020422323624837, 10010000010011111111010010100000100101011101001110111110000010000100001000010001001011011100011111011001011101001101101110000101";
	N_in <= "01010101110000000111010101011101010001000110111011111010000011111100100111001000110000010111011011001011001011101100101001000010";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10101011110111001011101111000000000000110010111110100111011101111000111010010100001101110000000010110000001110101000111100000001";
	wait for 33409 * clk_period;
	ASSERT(C_out = "10010000010011111111010010100000100101011101001110111110000010000100001000010001001011011100011111011001011101001101101110000101") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=191823984475670677583965020422323624837, exp=8940890154698342166679223776836487973, mod=228444100611487427329574816502404255489";
	REPORT "Expected output is 113983681069878420564395489959401671234, 01010101110000000111010101011101010001000110111011111010000011111100100111001000110000010111011011001011001011101100101001000010";
	N_in <= "10010000010011111111010010100000100101011101001110111110000010000100001000010001001011011100011111011001011101001101101110000101";
	Exp_in <= "00000110101110011111001111101011001101101111010010110101100000111100110010110011111110110110101000100011111011101000101100100101";
	M_in <= "10101011110111001011101111000000000000110010111110100111011101111000111010010100001101110000000010110000001110101000111100000001";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01010101110000000111010101011101010001000110111011111010000011111100100111001000110000010111011011001011001011101100101001000010") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=91501942807477730556433209096500104405, exp=65537, mod=237053248713799407909715617221250627043";
	REPORT "Expected output is 150892209896796217470381325386033495586, 01110001100001001100100001010100101000111100011111101011100001010011111000010011001001100111110011110101100101010111111000100010";
	N_in <= "01000100110101101010001000010110111010111110000110001000101101010011011001001101101001011100101011111100110010110100110011010101";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10110010010101101100101110000101110110101110110111010000011001001011100011110001101111001010110000110001001111111011010111100011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01110001100001001100100001010100101000111100011111101011100001010011111000010011001001100111110011110101100101010111111000100010") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=150892209896796217470381325386033495586, exp=159101335092011852019938343506938471793, mod=237053248713799407909715617221250627043";
	REPORT "Expected output is 91501942807477730556433209096500104405, 01000100110101101010001000010110111010111110000110001000101101010011011001001101101001011100101011111100110010110100110011010101";
	N_in <= "01110001100001001100100001010100101000111100011111101011100001010011111000010011001001100111110011110101100101010111111000100010";
	Exp_in <= "01110111101100011100110101110011100011111001011011100001101010001010101111111110011111111101011000010100010010001010010101110001";
	M_in <= "10110010010101101100101110000101110110101110110111010000011001001011100011110001101111001010110000110001001111111011010111100011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01000100110101101010001000010110111010111110000110001000101101010011011001001101101001011100101011111100110010110100110011010101") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=122431947429154588237871574947063942366, exp=65537, mod=171629935498219046480254733814521100511";
	REPORT "Expected output is 120187189805589358192985198612914536802, 01011010011010110011010111110101100010010011111001101000100100001011100010110010100111100101111000111111101110101000000101100010";
	N_in <= "01011100000110111000100100001110000001111110110000101100100101011001110101001001000101011001110110011011111101000100110011011110";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10000001000111101011100100100100011110110111110101110101101111101110110001001000011100010000101110100110000011110111100011011111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01011010011010110011010111110101100010010011111001101000100100001011100010110010100111100101111000111111101110101000000101100010") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=120187189805589358192985198612914536802, exp=137538071355584877117206977349970565561, mod=171629935498219046480254733814521100511";
	REPORT "Expected output is 122431947429154588237871574947063942366, 01011100000110111000100100001110000001111110110000101100100101011001110101001001000101011001110110011011111101000100110011011110";
	N_in <= "01011010011010110011010111110101100010010011111001101000100100001011100010110010100111100101111000111111101110101000000101100010";
	Exp_in <= "01100111011110001101111001110111100011001111101010111010011000110111000010011111111001001101110110001000011000000001100110111001";
	M_in <= "10000001000111101011100100100100011110110111110101110101101111101110110001001000011100010000101110100110000011110111100011011111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01011100000110111000100100001110000001111110110000101100100101011001110101001001000101011001110110011011111101000100110011011110") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=110245106113188858792990010842830825448, exp=65537, mod=230528543938941297765277192975286570351";
	REPORT "Expected output is 51817883121391364737874263430250102613, 00100110111110111100001011100010111110001111000110110011111010100101101110101111100010000101000111110001100011111111111101010101";
	N_in <= "01010010111100000110111101100011010001100011000100011000100111111100000110111110111101000110110011101000010101110110011111101000";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10101101011011100010111010111101100111011000001100000100100110010100001100110011110100000111010111110100101001001000110101101111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "00100110111110111100001011100010111110001111000110110011111010100101101110101111100010000101000111110001100011111111111101010101") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=51817883121391364737874263430250102613, exp=218881992998528482849611070024093421249, mod=230528543938941297765277192975286570351";
	REPORT "Expected output is 110245106113188858792990010842830825448, 01010010111100000110111101100011010001100011000100011000100111111100000110111110111101000110110011101000010101110110011111101000";
	N_in <= "00100110111110111100001011100010111110001111000110110011111010100101101110101111100010000101000111110001100011111111111101010101";
	Exp_in <= "10100100101010110010001101110010001000100110011001001110001000011011101010110110010100011001110011010010110111100100111011000001";
	M_in <= "10101101011011100010111010111101100111011000001100000100100110010100001100110011110100000111010111110100101001001000110101101111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01010010111100000110111101100011010001100011000100011000100111111100000110111110111101000110110011101000010101110110011111101000") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=128248564527951816691210905197506418122, exp=65537, mod=183626071149567297216181039737162798929";
	REPORT "Expected output is 159967332071542467689016557811837697627, 01111000010110001001011001100110001000111101010000010110100000011100100110010011001101100011100011010100110110111111111001011011";
	N_in <= "01100000011110111100011001101011010011110001110110101110001001110001000110000011011111001011001100000010100100110101010111001010";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10001010001001010001100001001011010110001111110011101011011011000011100011000111110001010111000101101010110100011001011101010001";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01111000010110001001011001100110001000111101010000010110100000011100100110010011001101100011100011010100110110111111111001011011") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=159967332071542467689016557811837697627, exp=105439924157354113268254690572630839297, mod=183626071149567297216181039737162798929";
	REPORT "Expected output is 128248564527951816691210905197506418122, 01100000011110111100011001101011010011110001110110101110001001110001000110000011011111001011001100000010100100110101010111001010";
	N_in <= "01111000010110001001011001100110001000111101010000010110100000011100100110010011001101100011100011010100110110111111111001011011";
	Exp_in <= "01001111010100101111110110100000010001100111100011110100101011111110101101000101111010110100110001100000100111010101000000000001";
	M_in <= "10001010001001010001100001001011010110001111110011101011011011000011100011000111110001010111000101101010110100011001011101010001";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01100000011110111100011001101011010011110001110110101110001001110001000110000011011111001011001100000010100100110101010111001010") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=141210003319477568027141702228654499670, exp=65537, mod=199073371188683318783368425487617891263";
	REPORT "Expected output is 73074949301072757149911567424758181154, 00110110111110011011100100101010011110010101011011001110000010001010000000001010110001101010111101001001110110110110110100100010";
	N_in <= "01101010001111000000111010110000101101111100010010000110101010101110011111101001111101111101001010001010011000010010011101010110";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10010101110001000010001011111100110100100010001101010001100101101000000000101100111001001100101010011100010001100001101110111111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "00110110111110011011100100101010011110010101011011001110000010001010000000001010110001101010111101001001110110110110110100100010") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=73074949301072757149911567424758181154, exp=80210132285706878705231396487593124833, mod=199073371188683318783368425487617891263";
	REPORT "Expected output is 141210003319477568027141702228654499670, 01101010001111000000111010110000101101111100010010000110101010101110011111101001111101111101001010001010011000010010011101010110";
	N_in <= "00110110111110011011100100101010011110010101011011001110000010001010000000001010110001101010111101001001110110110110110100100010";
	Exp_in <= "00111100010101111110100011011001000000010011101001100101110100100011101010111000001100100110001111110010011001101110001111100001";
	M_in <= "10010101110001000010001011111100110100100010001101010001100101101000000000101100111001001100101010011100010001100001101110111111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01101010001111000000111010110000101101111100010010000110101010101110011111101001111101111101001010001010011000010010011101010110") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=107401001106785305971232445883392932254, exp=65537, mod=223074455232137063705596207297494751693";
	REPORT "Expected output is 94841964166923530826419522747834381570, 01000111010110011110010111011011010010100110000000011011011110001010010110000010000110110001110101010010110001010011010100000010";
	N_in <= "01010000110011001010111000101111010001101001111100010010100110100100101100111110010101101001110111001011000011110011100110011110";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10100111110100101001001111001010111110100100110000010101111100100000001111110101101011010101101111000000011011111001100111001101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01000111010110011110010111011011010010100110000000011011011110001010010110000010000110110001110101010010110001010011010100000010") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=94841964166923530826419522747834381570, exp=3662482472950844259723435097945114497, mod=223074455232137063705596207297494751693";
	REPORT "Expected output is 107401001106785305971232445883392932254, 01010000110011001010111000101111010001101001111100010010100110100100101100111110010101101001110111001011000011110011100110011110";
	N_in <= "01000111010110011110010111011011010010100110000000011011011110001010010110000010000110110001110101010010110001010011010100000010";
	Exp_in <= "00000010110000010101111001010011110100101101000000110100111110111100100100110001000011101011011110000110101111011000011110000001";
	M_in <= "10100111110100101001001111001010111110100100110000010101111100100000001111110101101011010101101111000000011011111001100111001101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01010000110011001010111000101111010001101001111100010010100110100100101100111110010101101001110111001011000011110011100110011110") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=130315117460580382977070245191709535377, exp=65537, mod=297378603495393398829858271993873204387";
	REPORT "Expected output is 146388427224630179837896410739281075206, 01101110001000010110001010110011011011011100011111100111101110010001100010111110100110011010010001010001100001011001110000000110";
	N_in <= "01100010000010011100011101011000011000100000101010100010001010110111101101110101010111111101010000011110011010101010110010010001";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "11011111101110010000100100100101100011000011101101110010110011110001011001101101111010101110001101110000000011101000010010100011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01101110001000010110001010110011011011011100011111100111101110010001100010111110100110011010010001010001100001011001110000000110") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=146388427224630179837896410739281075206, exp=225821153854391309729346882542430915569, mod=297378603495393398829858271993873204387";
	REPORT "Expected output is 130315117460580382977070245191709535377, 01100010000010011100011101011000011000100000101010100010001010110111101101110101010111111101010000011110011010101010110010010001";
	N_in <= "01101110001000010110001010110011011011011100011111100111101110010001100010111110100110011010010001010001100001011001110000000110";
	Exp_in <= "10101001111000111001001001111101100011111110001011101000111111011100011000000000001001001000010000011010010001010000101111110001";
	M_in <= "11011111101110010000100100100101100011000011101101110010110011110001011001101101111010101110001101110000000011101000010010100011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01100010000010011100011101011000011000100000101010100010001010110111101101110101010111111101010000011110011010101010110010010001") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=114083607119984844524163149115957069507, exp=65537, mod=175917918563506049153379437745254583449";
	REPORT "Expected output is 29262888442581917127065487406442606025, 00010110000000111101001111001010101010001011110111010011000000000110010000110000101101110110101001110001000000011110110111001001";
	N_in <= "01010101110100111011010000011001010101100011100000000011010110110011100110001111010001001101010010110110001110100100011011000011";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10000100010110001000111100000111101110001011111010010010011100111000111100010000100011010100001100001101101010100100110010011001";
	wait for 33409 * clk_period;
	ASSERT(C_out = "00010110000000111101001111001010101010001011110111010011000000000110010000110000101101110110101001110001000000011110110111001001") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=29262888442581917127065487406442606025, exp=70550233510911843449935873972166067773, mod=175917918563506049153379437745254583449";
	REPORT "Expected output is 114083607119984844524163149115957069507, 01010101110100111011010000011001010101100011100000000011010110110011100110001111010001001101010010110110001110100100011011000011";
	N_in <= "00010110000000111101001111001010101010001011110111010011000000000110010000110000101101110110101001110001000000011110110111001001";
	Exp_in <= "00110101000100110111101100010001001000101011001100110010111011011111000000001010111010110001111001011111110000100000011000111101";
	M_in <= "10000100010110001000111100000111101110001011111010010010011100111000111100010000100011010100001100001101101010100100110010011001";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01010101110100111011010000011001010101100011100000000011010110110011100110001111010001001101010010110110001110100100011011000011") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=154722199386510637376774541998221403368, exp=65537, mod=206700370561945314919476792010479762097";
	REPORT "Expected output is 15782068964898419312304707877977096869, 00001011110111111000010000010011010110111100101011001101010010011110011011011111111110111010000000011110110101101000001010100101";
	N_in <= "01110100011001100110100101100100010000001101010110001101001111110101001110110100011101110011100100011000100110111010010011101000";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10011011100000010000101100010110111001010110111110111100000111011111110010000111001101001101111111100001100111111111101010110001";
	wait for 33409 * clk_period;
	ASSERT(C_out = "00001011110111111000010000010011010110111100101011001101010010011110011011011111111110111010000000011110110101101000001010100101") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=15782068964898419312304707877977096869, exp=193258238951786001114210143901440212673, mod=206700370561945314919476792010479762097";
	REPORT "Expected output is 154722199386510637376774541998221403368, 01110100011001100110100101100100010000001101010110001101001111110101001110110100011101110011100100011000100110111010010011101000";
	N_in <= "00001011110111111000010000010011010110111100101011001101010010011110011011011111111110111010000000011110110101101000001010100101";
	Exp_in <= "10010001011001000010111011010101001000101000000110111100110010000101011011011001000011010100111111101000001101101111111011000001";
	M_in <= "10011011100000010000101100010110111001010110111110111100000111011111110010000111001101001101111111100001100111111111101010110001";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01110100011001100110100101100100010000001101010110001101001111110101001110110100011101110011100100011000100110111010010011101000") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=147495708623944338425009786584638198039, exp=65537, mod=313646680610631121458743079196225278821";
	REPORT "Expected output is 183729479036049171972463008953371799599, 10001010001110010000001010110010010111101101111111001111100011000000111110110101000101001100000000010111000111010011000000101111";
	N_in <= "01101110111101101010001111100011100010100111000100101010000111010001001100100010100111110011001011101001001100001001000100010111";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "11101011111101100010011101000110001011010101010110101101111001000011101000101111110011010110010111100100100001011001001101100101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "10001010001110010000001010110010010111101101111111001111100011000000111110110101000101001100000000010111000111010011000000101111") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=183729479036049171972463008953371799599, exp=77525101533662107388192486420816272673, mod=313646680610631121458743079196225278821";
	REPORT "Expected output is 147495708623944338425009786584638198039, 01101110111101101010001111100011100010100111000100101010000111010001001100100010100111110011001011101001001100001001000100010111";
	N_in <= "10001010001110010000001010110010010111101101111111001111100011000000111110110101000101001100000000010111000111010011000000101111";
	Exp_in <= "00111010010100101100101010011100010111110000001001001001100010000100101011010101101110010110100110011111010001110001110100100001";
	M_in <= "11101011111101100010011101000110001011010101010110101101111001000011101000101111110011010110010111100100100001011001001101100101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01101110111101101010001111100011100010100111000100101010000111010001001100100010100111110011001011101001001100001001000100010111") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=132923046793359866552402336969101063382, exp=65537, mod=216951557236670656054676569872634358129";
	REPORT "Expected output is 59344469253135044347240703176317999304, 00101100101001010101010000111011110000100001101010010000000100000101011100101101010100111001001000001111110010100001100011001000";
	N_in <= "01100100000000000000110000110000010010100101001000101100111010101010111101011111110011010110000001110011001001101011010011010110";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10100011001101110101100110011101010010110001001001111010001101010101000110001011000110100000101100110011001100100010100101110001";
	wait for 33409 * clk_period;
	ASSERT(C_out = "00101100101001010101010000111011110000100001101010010000000100000101011100101101010100111001001000001111110010100001100011001000") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=59344469253135044347240703176317999304, exp=163191188444636668124173781100389953829, mod=216951557236670656054676569872634358129";
	REPORT "Expected output is 132923046793359866552402336969101063382, 01100100000000000000110000110000010010100101001000101100111010101010111101011111110011010110000001110011001001101011010011010110";
	N_in <= "00101100101001010101010000111011110000100001101010010000000100000101011100101101010100111001001000001111110010100001100011001000";
	Exp_in <= "01111010110001010111101011001010001111111001101100100001011110011001100000101110110001111111111011001111010110110111000100100101";
	M_in <= "10100011001101110101100110011101010010110001001001111010001101010101000110001011000110100000101100110011001100100010100101110001";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01100100000000000000110000110000010010100101001000101100111010101010111101011111110011010110000001110011001001101011010011010110") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=110474766028653274372647525965239121593, exp=65537, mod=289358127278560880418338415394372222319";
	REPORT "Expected output is 27855339526873030404738328524381990675, 00010100111101001011111001000101101010111010011101100101101110110011010010111001111110000101110101001000111000111010111100010011";
	N_in <= "01010011000111001010101001111110111011110110000111010011111110010010000100010001100000010110001101010110011110110111011010111001";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "11011001101100000101100100100011011111010000010011101111100101011010111001110011011001101011110010001111010111000111110101101111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "00010100111101001011111001000101101010111010011101100101101110110011010010111001111110000101110101001000111000111010111100010011") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=27855339526873030404738328524381990675, exp=118040031322647132622620632432866545353, mod=289358127278560880418338415394372222319";
	REPORT "Expected output is 110474766028653274372647525965239121593, 01010011000111001010101001111110111011110110000111010011111110010010000100010001100000010110001101010110011110110111011010111001";
	N_in <= "00010100111101001011111001000101101010111010011101100101101110110011010010111001111110000101110101001000111000111010111100010011";
	Exp_in <= "01011000110011011010111011011111011000100100110111010100001001001101001110111010000000111110101111000111100100001100111011001001";
	M_in <= "11011001101100000101100100100011011111010000010011101111100101011010111001110011011001101011110010001111010111000111110101101111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01010011000111001010101001111110111011110110000111010011111110010010000100010001100000010110001101010110011110110111011010111001") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=122111708942321626124448720633272088421, exp=65537, mod=245796187182256924961155953330036507889";
	REPORT "Expected output is 61942165735632647975335569205746037241, 00101110100110011010000010001110111011111101110111000110100111100100100000111111100010101101010100100110010010010111000111111001";
	N_in <= "01011011110111011101110000010100000100011011011010100001001111110001111100000110101100101100110011100110010000100011011101100101";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10111000111010101001111110101011100001110000100111101110110000000011001110101111010011011100001111001110010000011000010011110001";
	wait for 33409 * clk_period;
	ASSERT(C_out = "00101110100110011010000010001110111011111101110111000110100111100100100000111111100010101101010100100110010010010111000111111001") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=61942165735632647975335569205746037241, exp=21962898395399492668661998126608598913, mod=245796187182256924961155953330036507889";
	REPORT "Expected output is 122111708942321626124448720633272088421, 01011011110111011101110000010100000100011011011010100001001111110001111100000110101100101100110011100110010000100011011101100101";
	N_in <= "00101110100110011010000010001110111011111101110111000110100111100100100000111111100010101101010100100110010010010111000111111001";
	Exp_in <= "00010000100001011110011001111110100011010011001001110110000000011010111100100100100101001100101011110101111010101100011110000001";
	M_in <= "10111000111010101001111110101011100001110000100111101110110000000011001110101111010011011100001111001110010000011000010011110001";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01011011110111011101110000010100000100011011011010100001001111110001111100000110101100101100110011100110010000100011011101100101") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=107844471414724646263986568763593548763, exp=65537, mod=184262739251326738353309597355218499171";
	REPORT "Expected output is 10863739982750649923101813654205021994, 00001000001011000100011110111100000111000010110010000000001110111010000011011111001011011011010011101011010110001011111100101010";
	N_in <= "01010001001000100001011011110101011111100010100101101010011111011101000110111001100000000001111100111111111110010110001111011011";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10001010100111111011011001110100100011001000001101000100011110101010100100011101110010001001001001010101010101101111011001100011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "00001000001011000100011110111100000111000010110010000000001110111010000011011111001011011011010011101011010110001011111100101010") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=10863739982750649923101813654205021994, exp=45724780329345663408868247064506165921, mod=184262739251326738353309597355218499171";
	REPORT "Expected output is 107844471414724646263986568763593548763, 01010001001000100001011011110101011111100010100101101010011111011101000110111001100000000001111100111111111110010110001111011011";
	N_in <= "00001000001011000100011110111100000111000010110010000000001110111010000011011111001011011011010011101011010110001011111100101010";
	Exp_in <= "00100010011001100100010110111001101000000101000011000110110000000000011110001101001010100011100001011001111010100110101010100001";
	M_in <= "10001010100111111011011001110100100011001000001101000100011110101010100100011101110010001001001001010101010101101111011001100011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01010001001000100001011011110101011111100010100101101010011111011101000110111001100000000001111100111111111110010110001111011011") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=153211065691166335146442892894115225436, exp=65537, mod=229551668576583000904684805205753644501";
	REPORT "Expected output is 220046677895706813851531689748494677149, 10100101100010110111001011011000010000000011110110001001011111110000000000010010110110111110100000101011010010011111010010011101";
	N_in <= "01110011010000110110000010111111100010010100000100100001101010111000111001011011100110011110011001000011101100000101111101011100";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10101100101100100000101100010001000101111101001110000101011001100101100000001000010110100110010010010101011010001100010111010101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "10100101100010110111001011011000010000000011110110001001011111110000000000010010110110111110100000101011010010011111010010011101") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=220046677895706813851531689748494677149, exp=152938707245188521601402953639743236097, mod=229551668576583000904684805205753644501";
	REPORT "Expected output is 153211065691166335146442892894115225436, 01110011010000110110000010111111100010010100000100100001101010111000111001011011100110011110011001000011101100000101111101011100";
	N_in <= "10100101100010110111001011011000010000000011110110001001011111110000000000010010110110111110100000101011010010011111010010011101";
	Exp_in <= "01110011000011101110110001110000101001101111111100110110100010000110111001001011011100101000100001011111001111001010100000000001";
	M_in <= "10101100101100100000101100010001000101111101001110000101011001100101100000001000010110100110010010010101011010001100010111010101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01110011010000110110000010111111100010010100000100100001101010111000111001011011100110011110011001000011101100000101111101011100") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=140434737910795038188512766108771051826, exp=65537, mod=275214457394938630335103116379705415627";
	REPORT "Expected output is 214965929865586331908816366353781542238, 10100001101110001110111010100000011010000011011011100011010111001111011101101000111011011100111011011101010010101100110101011110";
	N_in <= "01101001101001101011111100100111100100001000011101010110011100011100001000111010001011101110011100001010010110000110100100110010";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "11001111000011000110000001011111110110010000001001111001001100010011011000001001111111011111110000110010011110011001011111001011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "10100001101110001110111010100000011010000011011011100011010111001111011101101000111011011100111011011101010010101100110101011110") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=214965929865586331908816366353781542238, exp=86654108798763425723988983058355672673, mod=275214457394938630335103116379705415627";
	REPORT "Expected output is 140434737910795038188512766108771051826, 01101001101001101011111100100111100100001000011101010110011100011100001000111010001011101110011100001010010110000110100100110010";
	N_in <= "10100001101110001110111010100000011010000011011011100011010111001111011101101000111011011100111011011101010010101100110101011110";
	Exp_in <= "01000001001100001111100101101011010101000110110111010101111011001000101100101101111101011001001101101100001101110101011001100001";
	M_in <= "11001111000011000110000001011111110110010000001001111001001100010011011000001001111111011111110000110010011110011001011111001011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01101001101001101011111100100111100100001000011101010110011100011100001000111010001011101110011100001010010110000110100100110010") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=108922376033674591478521157283659701450, exp=65537, mod=177003730340354578348766012138222195959";
	REPORT "Expected output is 30210489098733181888354784057426944020, 00010110101110100101010000011100011100010000100010101101101010010010001111000011101100001000101010001001111001111010000000010100";
	N_in <= "01010001111100011010111111000010100000100000101000101011011001110111010111000111010100110101011100010110101111001101110011001010";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10000101001010011010110110101111000110011100000101101110000010101001100101010001010010111001100010100011100011110001010011110111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "00010110101110100101010000011100011100010000100010101101101010010010001111000011101100001000101010001001111001111010000000010100") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=30210489098733181888354784057426944020, exp=163821021217397001571986237185000647425, mod=177003730340354578348766012138222195959";
	REPORT "Expected output is 108922376033674591478521157283659701450, 01010001111100011010111111000010100000100000101000101011011001110111010111000111010100110101011100010110101111001101110011001010";
	N_in <= "00010110101110100101010000011100011100010000100010101101101010010010001111000011101100001000101010001001111001111010000000010100";
	Exp_in <= "01111011001111101100011111110001011101111111010011111110110010011100001111111000010001001001011101100011111010101010101100000001";
	M_in <= "10000101001010011010110110101111000110011100000101101110000010101001100101010001010010111001100010100011100011110001010011110111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01010001111100011010111111000010100000100000101000101011011001110111010111000111010100110101011100010110101111001101110011001010") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=150173681022001669295078213130513050228, exp=65537, mod=207672510739458011785321106542614459157";
	REPORT "Expected output is 191703148539381144354797920412859526428, 10010000001110001010111011110100101001011101110101011000111110111011100000000100011000101101011000010110110011100110110100011100";
	N_in <= "01110000111110100110011000011111001110001110001001010011111100100011110011010011111101001111101000000010010111000110101001110100";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10011100001111000100010101001100111110111011001000011000101100110100101110110010111000101110011100011100000110101011001100010101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "10010000001110001010111011110100101001011101110101011000111110111011100000000100011000101101011000010110110011100110110100011100") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=191703148539381144354797920412859526428, exp=201914832603235798082782087861739902433, mod=207672510739458011785321106542614459157";
	REPORT "Expected output is 150173681022001669295078213130513050228, 01110000111110100110011000011111001110001110001001010011111100100011110011010011111101001111101000000010010111000110101001110100";
	N_in <= "10010000001110001010111011110100101001011101110101011000111110111011100000000100011000101101011000010110110011100110110100011100";
	Exp_in <= "10010111111001110110000111011001111111111011111010100001100010111000001100110001000100010100100100010101111011101101010111100001";
	M_in <= "10011100001111000100010101001100111110111011001000011000101100110100101110110010111000101110011100011100000110101011001100010101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01110000111110100110011000011111001110001110001001010011111100100011110011010011111101001111101000000010010111000110101001110100") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=148570955396077224098934017754928005333, exp=65537, mod=174342308227888794746656368580683901391";
	REPORT "Expected output is 165196274293581641506118484531514997973, 01111100010001111010010100100111101001110110101011010111011000111001000010110001111001110100110101110011100111000111110011010101";
	N_in <= "01101111110001011011100110100101110100000001001110110101111011001101110110011110011111100010110011111101101011000100000011010101";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10000011001010010001101101110001011001000011110111001111010111111110110100010001110010110101001010010011000011000010100111001111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01111100010001111010010100100111101001110110101011010111011000111001000010110001111001110100110101110011100111000111110011010101") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=165196274293581641506118484531514997973, exp=20225591184470428995358265017600246601, mod=174342308227888794746656368580683901391";
	REPORT "Expected output is 148570955396077224098934017754928005333, 01101111110001011011100110100101110100000001001110110101111011001101110110011110011111100010110011111101101011000100000011010101";
	N_in <= "01111100010001111010010100100111101001110110101011010111011000111001000010110001111001110100110101110011100111000111110011010101";
	Exp_in <= "00001111001101110100111010100010101110100000000101011101101100110101100111100000100011000001011010001000101011110000001101001001";
	M_in <= "10000011001010010001101101110001011001000011110111001111010111111110110100010001110010110101001010010011000011000010100111001111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01101111110001011011100110100101110100000001001110110101111011001101110110011110011111100010110011111101101011000100000011010101") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=109831774592829711927185006288292504876, exp=65537, mod=207513964353103747853255107762289226169";
	REPORT "Expected output is 200048749603740712371201535544966174478, 10010110011111111111110011011011001101100011100101111110101010110110010110110111111011110100101010000110001111101101011100001110";
	N_in <= "01010010101000001101010010010010000010011000101011110001010111101101110110011111001101110011001111111101010111110110010100101100";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10011100000111011011110001011100001111111101101110000001111010001100100101101011011000101101000010001010110001011011000110111001";
	wait for 33409 * clk_period;
	ASSERT(C_out = "10010110011111111111110011011011001101100011100101111110101010110110010110110111111011110100101010000110001111101101011100001110") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=200048749603740712371201535544966174478, exp=105794537085400650267436726233678238673, mod=207513964353103747853255107762289226169";
	REPORT "Expected output is 109831774592829711927185006288292504876, 01010010101000001101010010010010000010011000101011110001010111101101110110011111001101110011001111111101010111110110010100101100";
	N_in <= "10010110011111111111110011011011001101100011100101111110101010110110010110110111111011110100101010000110001111101101011100001110";
	Exp_in <= "01001111100101110100100101100100101011101001100110110110100001111111000111011011110010000111000111000110000010000101001111010001";
	M_in <= "10011100000111011011110001011100001111111101101110000001111010001100100101101011011000101101000010001010110001011011000110111001";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01010010101000001101010010010010000010011000101011110001010111101101110110011111001101110011001111111101010111110110010100101100") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=135526300806440520998262349569195207336, exp=65537, mod=172975787377627249077610378068618912997";
	REPORT "Expected output is 33947633491898638170759168152698329419, 00011001100010100001001110001110001011110011101001100100101101001010010111010101110111110111110110010111100001111001100101001011";
	N_in <= "01100101111101010110101010000101010111011110010101011011110101010001000001101001111111101000001111111011101100110110101010101000";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10000010001000011110110011000011011001000111101111111011000000100011010001110110001111011100100100110100011011000010010011100101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "00011001100010100001001110001110001011110011101001100100101101001010010111010101110111110111110110010111100001111001100101001011") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=33947633491898638170759168152698329419, exp=168026985916879105215551255777796568553, mod=172975787377627249077610378068618912997";
	REPORT "Expected output is 135526300806440520998262349569195207336, 01100101111101010110101010000101010111011110010101011011110101010001000001101001111111101000001111111011101100110110101010101000";
	N_in <= "00011001100010100001001110001110001011110011101001100100101101001010010111010101110111110111110110010111100001111001100101001011";
	Exp_in <= "01111110011010001101001000000011011001000010001100000011010000011001010101011111101101001110110110100011100011100011010111101001";
	M_in <= "10000010001000011110110011000011011001000111101111111011000000100011010001110110001111011100100100110100011011000010010011100101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01100101111101010110101010000101010111011110010101011011110101010001000001101001111111101000001111111011101100110110101010101000") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=99677357746016251962041102050411740407, exp=65537, mod=174606746752416730309072136455855708759";
	REPORT "Expected output is 134000035141197855047462146185264110950, 01100100110011110111011111010000010101101000111101000110101010010001111011001010111010000010011101110111101101000001110101100110";
	N_in <= "01001010111111010010100100101010100101011100000100000000010100100000010011100100100000101101100010000110111111001111110011110111";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10000011010111000000100101000100110100000001101101110010010101100100111010110100111101010000100011110010100101101001101001010111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01100100110011110111011111010000010101101000111101000110101010010001111011001010111010000010011101110111101101000001110101100110") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=134000035141197855047462146185264110950, exp=73924857746605841129073096540283860497, mod=174606746752416730309072136455855708759";
	REPORT "Expected output is 99677357746016251962041102050411740407, 01001010111111010010100100101010100101011100000100000000010100100000010011100100100000101101100010000110111111001111110011110111";
	N_in <= "01100100110011110111011111010000010101101000111101000110101010010001111011001010111010000010011101110111101101000001110101100110";
	Exp_in <= "00110111100111010110100011100011001101001000010011011010010011111111100000000001000010000110010000000111111100011111011000010001";
	M_in <= "10000011010111000000100101000100110100000001101101110010010101100100111010110100111101010000100011110010100101101001101001010111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01001010111111010010100100101010100101011100000100000000010100100000010011100100100000101101100010000110111111001111110011110111") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=167208775451516198672170269461213041433, exp=65537, mod=236163393091876799389320870257795287343";
	REPORT "Expected output is 37508440179887267062973264502484438690, 00011100001101111101110011100001001011100000001110111110110000000011111000101111011111010111111101011001001011010000111010100010";
	N_in <= "01111101110010110011110100011111011010101101001011010011011010110000001011001010110111111100101011010001111100110101001100011001";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10110001101010110110101001000000110111110101010000011101100001011000100001110110100110101101111101111011001101000100100100101111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "00011100001101111101110011100001001011100000001110111110110000000011111000101111011111010111111101011001001011010000111010100010") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=37508440179887267062973264502484438690, exp=24997565617564877176543869443532396161, mod=236163393091876799389320870257795287343";
	REPORT "Expected output is 167208775451516198672170269461213041433, 01111101110010110011110100011111011010101101001011010011011010110000001011001010110111111100101011010001111100110101001100011001";
	N_in <= "00011100001101111101110011100001001011100000001110111110110000000011111000101111011111010111111101011001001011010000111010100010";
	Exp_in <= "00010010110011100101101100100011110111001011111111010001100100101001111101000010001111001000001001110100110100000001011010000001";
	M_in <= "10110001101010110110101001000000110111110101010000011101100001011000100001110110100110101101111101111011001101000100100100101111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01111101110010110011110100011111011010101101001011010011011010110000001011001010110111111100101011010001111100110101001100011001") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=91739236726337134200328918152859262361, exp=65537, mod=210544450818395559485941271579284493737";
	REPORT "Expected output is 72735614352303821867832484239194509730, 00110110101110000101111010101001010001101011011101110111011101111001000010110011010000010001000000101100000110001101000110100010";
	N_in <= "01000101000001000101010110010101010000000110011011000011100100110101111000001110010111010100101001101100001110101001110110011001";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10011110011001010110001011100000111111010110000100111111011100101110001111110000110000100101101000100011010000000101010110101001";
	wait for 33409 * clk_period;
	ASSERT(C_out = "00110110101110000101111010101001010001101011011101110111011101111001000010110011010000010001000000101100000110001101000110100010") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=72735614352303821867832484239194509730, exp=166975110720449657308805500418776839773, mod=210544450818395559485941271579284493737";
	REPORT "Expected output is 91739236726337134200328918152859262361, 01000101000001000101010110010101010000000110011011000011100100110101111000001110010111010100101001101100001110101001110110011001";
	N_in <= "00110110101110000101111010101001010001101011011101110111011101111001000010110011010000010001000000101100000110001101000110100010";
	Exp_in <= "01111101100111100011110010001111111000001000001100101010011010101011100111101111101100011000010000010101100011110011011001011101";
	M_in <= "10011110011001010110001011100000111111010110000100111111011100101110001111110000110000100101101000100011010000000101010110101001";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01000101000001000101010110010101010000000110011011000011100100110101111000001110010111010100101001101100001110101001110110011001") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=143202895500040496005002920051609535161, exp=65537, mod=232404576723784748391049981915064102743";
	REPORT "Expected output is 226541647279369887722037693020635379047, 10101010011011100101010110001111000101101100100100011110100000010000111001001000100010010000111001011110111000111011010101100111";
	N_in <= "01101011101110111101111111011100011001000001001010110101001101010011101001010100100100101000011100100001110111011000001010111001";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10101110110101110111111001001100010110010110101101100010110001010111010000100001010000011110110011100001110100101110111101010111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "10101010011011100101010110001111000101101100100100011110100000010000111001001000100010010000111001011110111000111011010101100111") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=226541647279369887722037693020635379047, exp=223276765251074341210153933983872807825, mod=232404576723784748391049981915064102743";
	REPORT "Expected output is 143202895500040496005002920051609535161, 01101011101110111101111111011100011001000001001010110101001101010011101001010100100100101000011100100001110111011000001010111001";
	N_in <= "10101010011011100101010110001111000101101100100100011110100000010000111001001000100010010000111001011110111000111011010101100111";
	Exp_in <= "10100111111110011000101001110010011010011001101000111100110100001011000000010010110111010011011010101000110000010111001110010001";
	M_in <= "10101110110101110111111001001100010110010110101101100010110001010111010000100001010000011110110011100001110100101110111101010111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01101011101110111101111111011100011001000001001010110101001101010011101001010100100100101000011100100001110111011000001010111001") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=151135333693307530695101581201741915035, exp=65537, mod=205380933131878134586166284131985190681";
	REPORT "Expected output is 87423155427729966284559187176560198029, 01000001110001010001011001011000011100101010110000111000001110111000001110111011000010001100101100110001100000110000000110001101";
	N_in <= "01110001101100111001101101000010010111101111010001011101101000000101100000011000110111010011011001001000011010110010001110011011";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10011010100000101110110111001101001101010111001101011111001110101010111111101110111111101110010101010011011010101110111100011001";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01000001110001010001011001011000011100101010110000111000001110111000001110111011000010001100101100110001100000110000000110001101") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=87423155427729966284559187176560198029, exp=176230171882618473269046418115431685633, mod=205380933131878134586166284131985190681";
	REPORT "Expected output is 151135333693307530695101581201741915035, 01110001101100111001101101000010010111101111010001011101101000000101100000011000110111010011011001001000011010110010001110011011";
	N_in <= "01000001110001010001011001011000011100101010110000111000001110111000001110111011000010001100101100110001100000110000000110001101";
	Exp_in <= "10000100100101001011001001001110101100100111110110110011111111010000011011001011100011110101100110100101001001101101111000000001";
	M_in <= "10011010100000101110110111001101001101010111001101011111001110101010111111101110111111101110010101010011011010101110111100011001";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01110001101100111001101101000010010111101111010001011101101000000101100000011000110111010011011001001000011010110010001110011011") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=131083099394026673077449079289262796859, exp=65537, mod=188536688847263981303563932258335203351";
	REPORT "Expected output is 133913329738624987095797587376332031895, 01100100101111101100010011101000010011001110001101100100111011010010110101010000101001101101111000100100100101110100011110010111";
	N_in <= "01100010100111011010111111000111001001111000010001100100111011011100100110000101010101010101011110111110001100100111000000111011";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10001101110101101101100001110000100000001011011101100110101101111100000110001110010001110010011111101000111100000010000000010111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01100100101111101100010011101000010011001110001101100100111011010010110101010000101001101101111000100100100101110100011110010111") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=133913329738624987095797587376332031895, exp=137795731557671199969334439956268035217, mod=188536688847263981303563932258335203351";
	REPORT "Expected output is 131083099394026673077449079289262796859, 01100010100111011010111111000111001001111000010001100100111011011100100110000101010101010101011110111110001100100111000000111011";
	N_in <= "01100100101111101100010011101000010011001110001101100100111011010010110101010000101001101101111000100100100101110100011110010111";
	Exp_in <= "01100111101010100111111000011000100000111100101100000111100011100101101110000001001010010001001101110110111100011010110010010001";
	M_in <= "10001101110101101101100001110000100000001011011101100110101101111100000110001110010001110010011111101000111100000010000000010111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01100010100111011010111111000111001001111000010001100100111011011100100110000101010101010101011110111110001100100111000000111011") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=105608273409413658985169308893836586591, exp=65537, mod=181434525692383740295998533037515289071";
	REPORT "Expected output is 19140154612132413727807080450191175545, 00001110011001100100001001111011000110000010011101011001000010100101101001111101011101101000000101011011111010101010111101111001";
	N_in <= "01001111011100110110100111100010100100011011101001101010001101100101000100000100110010100010100110100110011101011010111001011111";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10001000011111110000010011000010110100010000111000000101000110011001101011010111010011000100111101111111010100110011000111101111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "00001110011001100100001001111011000110000010011101011001000010100101101001111101011101101000000101011011111010101010111101111001") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=19140154612132413727807080450191175545, exp=153191013918672723183767956626700770833, mod=181434525692383740295998533037515289071";
	REPORT "Expected output is 105608273409413658985169308893836586591, 01001111011100110110100111100010100100011011101001101010001101100101000100000100110010100010100110100110011101011010111001011111";
	N_in <= "00001110011001100100001001111011000110000010011101011001000010100101101001111101011101101000000101011011111010101010111101111001";
	Exp_in <= "01110011001111111000010000011110100101011111001100010111011101010000011111001011100100001101010111100111110001000001111000010001";
	M_in <= "10001000011111110000010011000010110100010000111000000101000110011001101011010111010011000100111101111111010100110011000111101111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01001111011100110110100111100010100100011011101001101010001101100101000100000100110010100010100110100110011101011010111001011111") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=124469930091882990953266069950118749420, exp=65537, mod=209925235847988879005662295672014606589";
	REPORT "Expected output is 116778402390958928037110947044692696971, 01010111110110101011001111000011100001101011110101011011100100101110001100100001000101101000010001110111001111011001111110001011";
	N_in <= "01011101101001000000100101011011100110011110110001001110000000100001010001101000001011011001110001111010001111111110010011101100";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10011101111011100010000100111001010001101100011000111110101101110011001111000000100100100010100011111011000010011001000011111101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01010111110110101011001111000011100001101011110101011011100100101110001100100001000101101000010001110111001111011001111110001011") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=116778402390958928037110947044692696971, exp=157079567889124107376830968935766892101, mod=209925235847988879005662295672014606589";
	REPORT "Expected output is 124469930091882990953266069950118749420, 01011101101001000000100101011011100110011110110001001110000000100001010001101000001011011001110001111010001111111110010011101100";
	N_in <= "01010111110110101011001111000011100001101011110101011011100100101110001100100001000101101000010001110111001111011001111110001011";
	Exp_in <= "01110110001011000110110010100001110111100010101010010011010100101110001000011111010110001011111101110111100001010001111001000101";
	M_in <= "10011101111011100010000100111001010001101100011000111110101101110011001111000000100100100010100011111011000010011001000011111101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01011101101001000000100101011011100110011110110001001110000000100001010001101000001011011001110001111010001111111110010011101100") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=149176772362218874633993551409003276355, exp=65537, mod=170710691922558067341512918363362509679";
	REPORT "Expected output is 27245876545453801588120428194147267397, 00010100011111110101110101101101010111001110110010100101001010011110111111001101110111001000110011001110011001101111001101000101";
	N_in <= "01110000001110100110011010111010111100000000111111000111001010001000010001111000010011111001010100101110001111101010100001000011";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10000000011011011010111011101111010111111111110011000110100110010110111100000010111011111001011100101001000100110100001101101111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "00010100011111110101110101101101010111001110110010100101001010011110111111001101110111001000110011001110011001101111001101000101") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=27245876545453801588120428194147267397, exp=133912700790983875277346620345504947073, mod=170710691922558067341512918363362509679";
	REPORT "Expected output is 149176772362218874633993551409003276355, 01110000001110100110011010111010111100000000111111000111001010001000010001111000010011111001010100101110001111101010100001000011";
	N_in <= "00010100011111110101110101101101010111001110110010100101001010011110111111001101110111001000110011001110011001101111001101000101";
	Exp_in <= "01100100101111101010010111100101110111010111010001011011000001111101010010100011001110001111001001011000110100101101101110000001";
	M_in <= "10000000011011011010111011101111010111111111110011000110100110010110111100000010111011111001011100101001000100110100001101101111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01110000001110100110011010111010111100000000111111000111001010001000010001111000010011111001010100101110001111101010100001000011") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=165670569628412269280971573671021621864, exp=65537, mod=257028066483625303712679302390526238061";
	REPORT "Expected output is 99953766894251456993065509139548391384, 01001011001100100110010100110000100001001110100101110101011100100111001010011000000000111000110010000011001101101100011111011000";
	N_in <= "01111100101000101111110110111000011010001010011100010101010110100100000000101010001000011000000110101101110111011011001001101000";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "11000001010111011100111000010011000110000111110110000000001011010001010010011000011011000110010100101000111000111101110101101101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01001011001100100110010100110000100001001110100101110101011100100111001010011000000000111000110010000011001101101100011111011000") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=99953766894251456993065509139548391384, exp=139022703216679887028476160677164368673, mod=257028066483625303712679302390526238061";
	REPORT "Expected output is 165670569628412269280971573671021621864, 01111100101000101111110110111000011010001010011100010101010110100100000000101010001000011000000110101101110111011011001001101000";
	N_in <= "01001011001100100110010100110000100001001110100101110101011100100111001010011000000000111000110010000011001101101100011111011000";
	Exp_in <= "01101000100101101100110001111000000101111010111100001010001101010011100000101101000000100101010100100100101101000100001100100001";
	M_in <= "11000001010111011100111000010011000110000111110110000000001011010001010010011000011011000110010100101000111000111101110101101101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01111100101000101111110110111000011010001010011100010101010110100100000000101010001000011000000110101101110111011011001001101000") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=152630371931377026717620176410579647167, exp=65537, mod=196060243432949451840762357818665775681";
	REPORT "Expected output is 47356199762405082096616964783155908283, 00100011101000000111100011101001110011000110000111000111100010011100010011011111101110110001110110101100101011110000111010111011";
	N_in <= "01110010110100111000101001010101110110110010100011100100000000101100000001110110000110000111010111011011000000010011101010111111";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10010011011111111101010001010001110011000100001011011001010111101000111111100100000110010001101000100110010100001011001001000001";
	wait for 33409 * clk_period;
	ASSERT(C_out = "00100011101000000111100011101001110011000110000111000111100010011100010011011111101110110001110110101100101011110000111010111011") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=47356199762405082096616964783155908283, exp=121952421129197009241660594567651177473, mod=196060243432949451840762357818665775681";
	REPORT "Expected output is 152630371931377026717620176410579647167, 01110010110100111000101001010101110110110010100011100100000000101100000001110110000110000111010111011011000000010011101010111111";
	N_in <= "00100011101000000111100011101001110011000110000111000111100010011100010011011111101110110001110110101100101011110000111010111011";
	Exp_in <= "01011011101111110010111010010101001101101100010111111010001000011001100000010110010100011110000011010111001010101011010000000001";
	M_in <= "10010011011111111101010001010001110011000100001011011001010111101000111111100100000110010001101000100110010100001011001001000001";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01110010110100111000101001010101110110110010100011100100000000101100000001110110000110000111010111011011000000010011101010111111") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=128800475760721843518907485429272260144, exp=65537, mod=210830533418527815966922892882026095737";
	REPORT "Expected output is 102101656307585970940500817846507115513, 01001100110100000001000001010000010011110101001110101010010011110101110011100110100101100011101011011100101010111001001111111001";
	N_in <= "01100000111001100001000110111110011011001000101101001001101001111100000111010110010010100100000101011000110101011010111000110000";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10011110100111000111101111010111000011010110001101101001000111111010000101011010101001111110110110100000100111101110010001111001";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01001100110100000001000001010000010011110101001110101010010011110101110011100110100101100011101011011100101010111001001111111001") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=102101656307585970940500817846507115513, exp=176273846509120522171162660379118046733, mod=210830533418527815966922892882026095737";
	REPORT "Expected output is 128800475760721843518907485429272260144, 01100000111001100001000110111110011011001000101101001001101001111100000111010110010010100100000101011000110101011010111000110000";
	N_in <= "01001100110100000001000001010000010011110101001110101010010011110101110011100110100101100011101011011100101010111001001111111001";
	Exp_in <= "10000100100111010001101110100001111110111100110010110001010011010101111110110000111101110111111111000110011010001000111000001101";
	M_in <= "10011110100111000111101111010111000011010110001101101001000111111010000101011010101001111110110110100000100111101110010001111001";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01100000111001100001000110111110011011001000101101001001101001111100000111010110010010100100000101011000110101011010111000110000") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=169482918641750193266520805340069216881, exp=65537, mod=204483075463039489635706770745022218499";
	REPORT "Expected output is 6050324858093110445349236835911232819, 00000100100011010100000000001011111010010011011001000100111100110111000110010011110110111001111011111001100011000110110100110011";
	N_in <= "01111111100000010011100100001001111010000101110111100000110001111000000011111000001001111001111101100110011110111100001001110001";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10011001110101100000001000000000001100011100001111111100111110100001010001011101011100010110111111001110010111000000000100000011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "00000100100011010100000000001011111010010011011001000100111100110111000110010011110110111001111011111001100011000110110100110011") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=6050324858093110445349236835911232819, exp=121634621875446411289733479016707589825, mod=204483075463039489635706770745022218499";
	REPORT "Expected output is 169482918641750193266520805340069216881, 01111111100000010011100100001001111010000101110111100000110001111000000011111000001001111001111101100110011110111100001001110001";
	N_in <= "00000100100011010100000000001011111010010011011001000100111100110111000110010011110110111001111011111001100011000110110100110011";
	Exp_in <= "01011011100000011111100111011110101100111011101110101001100100011111011011010100001100011000000010101001110100110000011011000001";
	M_in <= "10011001110101100000001000000000001100011100001111111100111110100001010001011101011100010110111111001110010111000000000100000011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01111111100000010011100100001001111010000101110111100000110001111000000011111000001001111001111101100110011110111100001001110001") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=114272429068568200083322727137624323421, exp=65537, mod=289950650526298553088093497097561371887";
	REPORT "Expected output is 141270909851944448028586107827372538208, 01101010010001111100100110011101001111000011011011110101111100010100010000011001101110111011110011000001100011011011100101100000";
	N_in <= "01010101111110000001000110111101011000111010110010100110010000101110011100101110100011100010110001110111111001011111010101011101";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "11011010001000100111011011001010010011000010110001111110010010101001111100011111111000000000000101110011101011001111010011101111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01101010010001111100100110011101001111000011011011110101111100010100010000011001101110111011110011000001100011011011100101100000") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=141270909851944448028586107827372538208, exp=194568712465409734289482667523568416337, mod=289950650526298553088093497097561371887";
	REPORT "Expected output is 114272429068568200083322727137624323421, 01010101111110000001000110111101011000111010110010100110010000101110011100101110100011100010110001110111111001011111010101011101";
	N_in <= "01101010010001111100100110011101001111000011011011110101111100010100010000011001101110111011110011000001100011011011100101100000";
	Exp_in <= "10010010011000001001001000101010010010100101011110001001000101100110001001000101110101111100110000010110100011011011011001010001";
	M_in <= "11011010001000100111011011001010010011000010110001111110010010101001111100011111111000000000000101110011101011001111010011101111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01010101111110000001000110111101011000111010110010100110010000101110011100101110100011100010110001110111111001011111010101011101") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=91977357235172032013093587542486682039, exp=65537, mod=235957421680162956462555042630296701093";
	REPORT "Expected output is 48864485689297448836793806065510882361, 00100100110000101111010100100110100111111101000110110111111011101000011100100101100111001000010011010110111000111001110000111001";
	N_in <= "01000101001100100011000111010100100111010010111001000000110111010110100100100000101010000101000101111001011001100000100110110111";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10110001100000111011111100010100001010011110011000111111001100101010101010011100011110011110110110110100000000001000100010100101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "00100100110000101111010100100110100111111101000110110111111011101000011100100101100111001000010011010110111000111001110000111001") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=48864485689297448836793806065510882361, exp=230344445492675368344934178242947143105, mod=235957421680162956462555042630296701093";
	REPORT "Expected output is 91977357235172032013093587542486682039, 01000101001100100011000111010100100111010010111001000000110111010110100100100000101010000101000101111001011001100000100110110111";
	N_in <= "00100100110000101111010100100110100111111101000110110111111011101000011100100101100111001000010011010110111000111001110000111001";
	Exp_in <= "10101101010010101011100111111100100010110011001010110100101100000100111011010111110001011010000100101111001000110101010111000001";
	M_in <= "10110001100000111011111100010100001010011110011000111111001100101010101010011100011110011110110110110100000000001000100010100101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01000101001100100011000111010100100111010010111001000000110111010110100100100000101010000101000101111001011001100000100110110111") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=134396470369257450997620053122546901505, exp=65537, mod=184576450819436289001524472161766668941";
	REPORT "Expected output is 137602762369047902174186361175707263716, 01100111100001010101001111111010111011110000100110111111110100101000111010100001011000111000110000100010101011001010001011100100";
	N_in <= "01100101000110111101000110010100011000100100111100110110001110011110011011000101010100101100011001100101111110111010001000000001";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10001010110111000010000110100001001101101110010100011000101100011101110100000101110101110000111111100110101100101111101010001101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01100111100001010101001111111010111011110000100110111111110100101000111010100001011000111000110000100010101011001010001011100100") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=137602762369047902174186361175707263716, exp=113153303699780151312046709129901250205, mod=184576450819436289001524472161766668941";
	REPORT "Expected output is 134396470369257450997620053122546901505, 01100101000110111101000110010100011000100100111100110110001110011110011011000101010100101100011001100101111110111010001000000001";
	N_in <= "01100111100001010101001111111010111011110000100110111111110100101000111010100001011000111000110000100010101011001010001011100100";
	Exp_in <= "01010101001000001000100010011001010111011001111011101011000101000011000100110110110111011111111011011101110010000001011010011101";
	M_in <= "10001010110111000010000110100001001101101110010100011000101100011101110100000101110101110000111111100110101100101111101010001101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01100101000110111101000110010100011000100100111100110110001110011110011011000101010100101100011001100101111110111010001000000001") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=143382123557734254678950589325996174662, exp=65537, mod=172810761380193137401959583259583989143";
	REPORT "Expected output is 157102307639601297272745442776265703454, 01110110001100001100110111001001110111101100001110011001101101010111001010101000011001100100111101011010100100101100000000011110";
	N_in <= "01101011110111100110010001111100100001000010100010000101010000010101000111111000000011100101010111111010110111111010110101000110";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10000010000000100010010001011010011110000000111101000001111101000011111111010100010100010111110001010000001011100100010110010111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01110110001100001100110111001001110111101100001110011001101101010111001010101000011001100100111101011010100100101100000000011110") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=157102307639601297272745442776265703454, exp=23111926446089885829817660089922735073, mod=172810761380193137401959583259583989143";
	REPORT "Expected output is 143382123557734254678950589325996174662, 01101011110111100110010001111100100001000010100010000101010000010101000111111000000011100101010111111010110111111010110101000110";
	N_in <= "01110110001100001100110111001001110111101100001110011001101101010111001010101000011001100100111101011010100100101100000000011110";
	Exp_in <= "00010001011000110011000111110011011110111000110100100110110101101001100011111001010011000010011101011101110011111100101111100001";
	M_in <= "10000010000000100010010001011010011110000000111101000001111101000011111111010100010100010111110001010000001011100100010110010111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01101011110111100110010001111100100001000010100010000101010000010101000111111000000011100101010111111010110111111010110101000110") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=136345945714578895352084234002766777115, exp=65537, mod=195213603457058976599229077284120815323";
	REPORT "Expected output is 136454551717013620196568138950149760469, 01100110101010000011000011010011000001100011000000011110111000010111110110010110110001100011001101111011110011010110010111010101";
	N_in <= "01100110100100110100011000100010100011011100101100111010101101000111100100001111110010010100000101100001110011000100101100011011";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10010010110111001100010110111110111101000001010111100010100111001110010111010110100000110010100001010001000111011110011011011011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01100110101010000011000011010011000001100011000000011110111000010111110110010110110001100011001101111011110011010110010111010101") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=136454551717013620196568138950149760469, exp=74672472421151585809074308833058331713, mod=195213603457058976599229077284120815323";
	REPORT "Expected output is 136345945714578895352084234002766777115, 01100110100100110100011000100010100011011100101100111010101101000111100100001111110010010100000101100001110011000100101100011011";
	N_in <= "01100110101010000011000011010011000001100011000000011110111000010111110110010110110001100011001101111011110011010110010111010101";
	Exp_in <= "00111000001011010110010100100011000001110010000100111011111110101011010111100110110101110111110010100011110000011001110001000001";
	M_in <= "10010010110111001100010110111110111101000001010111100010100111001110010111010110100000110010100001010001000111011110011011011011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01100110100100110100011000100010100011011100101100111010101101000111100100001111110010010100000101100001110011000100101100011011") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=134317519886564928539432497938359743256, exp=65537, mod=286717881484536854187231839071735398007";
	REPORT "Expected output is 13970961228362708440063659438216846444, 00001010100000101011010110010001111100010100111110101010010001011110100101101011111010000100000111101001111001000001110001101100";
	N_in <= "01100101000011001001110100000101001100100011010001000000111111101001000001111111110001100001100100110101100100010111001100011000";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "11010111101100111101101011111000011111101011110110010110010000001011000011000100110001100111000000110011101001000011111001110111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "00001010100000101011010110010001111100010100111110101010010001011110100101101011111010000100000111101001111001000001110001101100") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=13970961228362708440063659438216846444, exp=112544326124017128757606784484867465473, mod=286717881484536854187231839071735398007";
	REPORT "Expected output is 134317519886564928539432497938359743256, 01100101000011001001110100000101001100100011010001000000111111101001000001111111110001100001100100110101100100010111001100011000";
	N_in <= "00001010100000101011010110010001111100010100111110101010010001011110100101101011111010000100000111101001111001000001110001101100";
	Exp_in <= "01010100101010110011111110101111101111010010100000110100000101011111110101010110100111010100100100000111011100100110000100000001";
	M_in <= "11010111101100111101101011111000011111101011110110010110010000001011000011000100110001100111000000110011101001000011111001110111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01100101000011001001110100000101001100100011010001000000111111101001000001111111110001100001100100110101100100010111001100011000") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=132661752808201312184286541636668566249, exp=65537, mod=257368969124391078306549888792044614691";
	REPORT "Expected output is 23521800128361777458418762430651731087, 00010001101100100010001001001000101010101100000000101110000110010000010010001011001100001000111001111001110011101000110010001111";
	N_in <= "01100011110011011011100101100110100010010010011001001100111111001100000001110101101101100101111011111110110111010010101011101001";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "11000001100111110111010111011111010110010010011100010100001100000010100011111110001000111000011011010101000100011011010000100011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "00010001101100100010001001001000101010101100000000101110000110010000010010001011001100001000111001111001110011101000110010001111") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=23521800128361777458418762430651731087, exp=59169297615044942144140423953611040017, mod=257368969124391078306549888792044614691";
	REPORT "Expected output is 132661752808201312184286541636668566249, 01100011110011011011100101100110100010010010011001001100111111001100000001110101101101100101111011111110110111010010101011101001";
	N_in <= "00010001101100100010001001001000101010101100000000101110000110010000010010001011001100001000111001111001110011101000110010001111";
	Exp_in <= "00101100100000111001011110011010110110001010100101000110010101001111100110100001001010000011011000011101111100010010010100010001";
	M_in <= "11000001100111110111010111011111010110010010011100010100001100000010100011111110001000111000011011010101000100011011010000100011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01100011110011011011100101100110100010010010011001001100111111001100000001110101101101100101111011111110110111010010101011101001") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=92094543360962544252279523520596148073, exp=65537, mod=192720295454947370185957410183733506377";
	REPORT "Expected output is 179677576147531126038136996120782293604, 10000111001011001010010001110101111000011110111000010010001111111111100101111111010101111101110110010001011011011100101001100100";
	N_in <= "01000101010010001100001110001101011101110110000001011101100011011110111000101001110101000110001000010011111011111111111101101001";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10010000111111001001010000101011101000011111111111010111010010110110010100110011100101110110101011001111010010101111000101001001";
	wait for 33409 * clk_period;
	ASSERT(C_out = "10000111001011001010010001110101111000011110111000010010001111111111100101111111010101111101110110010001011011011100101001100100") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=179677576147531126038136996120782293604, exp=63679417704150102949765445081639732813, mod=192720295454947370185957410183733506377";
	REPORT "Expected output is 92094543360962544252279523520596148073, 01000101010010001100001110001101011101110110000001011101100011011110111000101001110101000110001000010011111011111111111101101001";
	N_in <= "10000111001011001010010001110101111000011110111000010010001111111111100101111111010101111101110110010001011011011100101001100100";
	Exp_in <= "00101111111010000011010110110001100000010011001011111111010101100010000001111000110011101101001111011001101010001100011001001101";
	M_in <= "10010000111111001001010000101011101000011111111111010111010010110110010100110011100101110110101011001111010010101111000101001001";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01000101010010001100001110001101011101110110000001011101100011011110111000101001110101000110001000010011111011111111111101101001") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=109127058252370095555465907379805189563, exp=65537, mod=171886624152636585929295642340878946921";
	REPORT "Expected output is 109084301535238047694412456892253071399, 01010010000100001101111101001101101010111111110101100010101100000010101000001110011000110111000100100010010111111110100000100111";
	N_in <= "01010010000110010001101101011111010100000010100101101101111011000000101000111010000001100111010000110100101100010111010110111011";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10000001010100000010100011011110110010100111100111111001000000000011000110111000111100100000111001101110001010111001001001101001";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01010010000100001101111101001101101010111111110101100010101100000010101000001110011000110111000100100010010111111110100000100111") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=109084301535238047694412456892253071399, exp=142800418469545511373247734805795063985, mod=171886624152636585929295642340878946921";
	REPORT "Expected output is 109127058252370095555465907379805189563, 01010010000110010001101101011111010100000010100101101101111011000000101000111010000001100111010000110100101100010111010110111011";
	N_in <= "01010010000100001101111101001101101010111111110101100010101100000010101000001110011000110111000100100010010111111110100000100111";
	Exp_in <= "01101011011011100101110000110110000100111100001101010111110001010111000011000100100110110100110111011000111111100100100010110001";
	M_in <= "10000001010100000010100011011110110010100111100111111001000000000011000110111000111100100000111001101110001010111001001001101001";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01010010000110010001101101011111010100000010100101101101111011000000101000111010000001100111010000110100101100010111010110111011") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=92106282370968335120447520903794720775, exp=65537, mod=231956804162469220138249298516206890923";
	REPORT "Expected output is 47506374572675868488149498024090573783, 00100011101111010110010100011010011000101111111110011010011011100100011001001001001100011001101001111100101010101001101111010111";
	N_in <= "01000101010010110000011001010100100110100110111110111000101111101001011111010001000111101000011101110110011111110000000000000111";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10101110100000010100000101101000000011110111100111111000000100011100111000111111110011001110110101001111111100110010111110101011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "00100011101111010110010100011010011000101111111110011010011011100100011001001001001100011001101001111100101010101001101111010111") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=47506374572675868488149498024090573783, exp=20078596060449637370355864076248281753, mod=231956804162469220138249298516206890923";
	REPORT "Expected output is 92106282370968335120447520903794720775, 01000101010010110000011001010100100110100110111110111000101111101001011111010001000111101000011101110110011111110000000000000111";
	N_in <= "00100011101111010110010100011010011000101111111110011010011011100100011001001001001100011001101001111100101010101001101111010111";
	Exp_in <= "00001111000110101111111100110111011010111100011110001010000100010111101000101101010010000011011110010000110000011111001010011001";
	M_in <= "10101110100000010100000101101000000011110111100111111000000100011100111000111111110011001110110101001111111100110010111110101011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01000101010010110000011001010100100110100110111110111000101111101001011111010001000111101000011101110110011111110000000000000111") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=126280015550946940280351265710884118649, exp=65537, mod=185204573713905628758585841890686924429";
	REPORT "Expected output is 129049999810114939417467963792847385034, 01100001000101100010000000111010101101000010001011111011000100000010000001111111100011011010001111011001001011011011000111001010";
	N_in <= "01011111000000001010010101110110000011111011111000100110100011110100001011100100011011111101101100111001111001011110000001111001";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10001011010101010001101001111010101111001000001011010011010111111111101101110111001101101111100111010000100001111111011010001101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01100001000101100010000000111010101101000010001011111011000100000010000001111111100011011010001111011001001011011011000111001010") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=129049999810114939417467963792847385034, exp=31970022161914862985031754560414042589, mod=185204573713905628758585841890686924429";
	REPORT "Expected output is 126280015550946940280351265710884118649, 01011111000000001010010101110110000011111011111000100110100011110100001011100100011011111101101100111001111001011110000001111001";
	N_in <= "01100001000101100010000000111010101101000010001011111011000100000010000001111111100011011010001111011001001011011011000111001010";
	Exp_in <= "00011000000011010011001111001001111101100001101010011011010000100001111001110110111000011100100110100101111111100100100111011101";
	M_in <= "10001011010101010001101001111010101111001000001011010011010111111111101101110111001101101111100111010000100001111111011010001101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01011111000000001010010101110110000011111011111000100110100011110100001011100100011011111101101100111001111001011110000001111001") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=99337639429939004548525630466393322883, exp=65537, mod=185835992198566931950671130854662988911";
	REPORT "Expected output is 10169996432107293027392445480368448831, 00000111101001101010101110001001011101101110010010011101110101111111001011001000011010010011010100001010101111011010010100111111";
	N_in <= "01001010101110111011101111000010100111001000110010111101100111000100111000001111000000101000011110110000000011110011010110000011";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10001011110011101011010111010000011101000101101001000100010101111111000110010001010111111010000000010000111101011110010001101111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "00000111101001101010101110001001011101101110010010011101110101111111001011001000011010010011010100001010101111011010010100111111") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=10169996432107293027392445480368448831, exp=24760362602467101763100549293599019937, mod=185835992198566931950671130854662988911";
	REPORT "Expected output is 99337639429939004548525630466393322883, 01001010101110111011101111000010100111001000110010111101100111000100111000001111000000101000011110110000000011110011010110000011";
	N_in <= "00000111101001101010101110001001011101101110010010011101110101111111001011001000011010010011010100001010101111011010010100111111";
	Exp_in <= "00010010101000001010110000100000111001100001111111010000110100100000111110111010010100101011011000111110100011101101001110100001";
	M_in <= "10001011110011101011010111010000011101000101101001000100010101111111000110010001010111111010000000010000111101011110010001101111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01001010101110111011101111000010100111001000110010111101100111000100111000001111000000101000011110110000000011110011010110000011") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=137229883547002831986236346442179540682, exp=65537, mod=229126654758483632321370712260190367117";
	REPORT "Expected output is 73843978820944862478186041931981569654, 00110111100011011101010100111111101001010001110111111001010000101010101110101011101101011001110001000000100011101011111001110110";
	N_in <= "01100111001111011000001110100010100010000011111001110100111011011000000001010001001110111001001001011100100100011111011011001010";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10101100011000000011000001000100100001110101010010010101100101010011000011011111010111011111000111011000111010110110110110001101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "00110111100011011101010100111111101001010001110111111001010000101010101110101011101101011001110001000000100011101011111001110110") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=73843978820944862478186041931981569654, exp=193833101806915933423011168480872619833, mod=229126654758483632321370712260190367117";
	REPORT "Expected output is 137229883547002831986236346442179540682, 01100111001111011000001110100010100010000011111001110100111011011000000001010001001110111001001001011100100100011111011011001010";
	N_in <= "00110111100011011101010100111111101001010001110111111001010000101010101110101011101101011001110001000000100011101011111001110110";
	Exp_in <= "10010001110100101110010111000010011100111000001000011000111001010010101001100100000110111100100010101101011100111101111100111001";
	M_in <= "10101100011000000011000001000100100001110101010010010101100101010011000011011111010111011111000111011000111010110110110110001101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01100111001111011000001110100010100010000011111001110100111011011000000001010001001110111001001001011100100100011111011011001010") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=111498348975957716648988340996667081735, exp=65537, mod=201127694995540430520877107238807323391";
	REPORT "Expected output is 65380972895495748854323751556393928614, 00110001001011111110101011010111011001101011000100010010101100000100000101100011110110111000011010001100011011110000011110100110";
	N_in <= "01010011111000011100110100001000000011111010011111110011001101010010101010100100101111110010111000111000111011000000010000000111";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10010111010011111100100011111000101000001000110110100110111100000101010001000100110101000011001110111110111010001100001011111111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "00110001001011111110101011010111011001101011000100010010101100000100000101100011110110111000011010001100011011110000011110100110") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=65380972895495748854323751556393928614, exp=70075679196914265013855683550736298577, mod=201127694995540430520877107238807323391";
	REPORT "Expected output is 111498348975957716648988340996667081735, 01010011111000011100110100001000000011111010011111110011001101010010101010100100101111110010111000111000111011000000010000000111";
	N_in <= "00110001001011111110101011010111011001101011000100010010101100000100000101100011110110111000011010001100011011110000011110100110";
	Exp_in <= "00110100101110000001010110111011100110101010010100000000000010111001100101111110001100100100001100000111011111000011001001010001";
	M_in <= "10010111010011111100100011111000101000001000110110100110111100000101010001000100110101000011001110111110111010001100001011111111";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01010011111000011100110100001000000011111010011111110011001101010010101010100100101111110010111000111000111011000000010000000111") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=162000219790812923746766626330535885843, exp=65537, mod=204469999776634988411550689937839242261";
	REPORT "Expected output is 151826681190665548186724815819402609618, 01110010001110001100000101010010100100101000001111111001001010110110101010000100110000011001000110011001001110111000001111010010";
	N_in <= "01111001111000000001101110000000011110111010000111000000010010011000011011011101011101111011100011001011010101010111110000010011";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10011001110100110111110101010001110101000101001001011100100100000000000010111011100111111111101101010111010101100011110000010101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01110010001110001100000101010010100100101000001111111001001010110110101010000100110000011001000110011001001110111000001111010010") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=151826681190665548186724815819402609618, exp=137906570794006740448448948353706885177, mod=204469999776634988411550689937839242261";
	REPORT "Expected output is 162000219790812923746766626330535885843, 01111001111000000001101110000000011110111010000111000000010010011000011011011101011101111011100011001011010101010111110000010011";
	N_in <= "01110010001110001100000101010010100100101000001111111001001010110110101010000100110000011001000110011001001110111000001111010010";
	Exp_in <= "01100111101111111101011011100100010111000001100111111000110000001100111000011001100111011000001001110100101100100000000000111001";
	M_in <= "10011001110100110111110101010001110101000101001001011100100100000000000010111011100111111111101101010111010101100011110000010101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01111001111000000001101110000000011110111010000111000000010010011000011011011101011101111011100011001011010101010111110000010011") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=141453349230748878185067692217169657844, exp=65537, mod=184822667877625730707730917278973060021";
	REPORT "Expected output is 169619234061427452515943317301574317356, 01111111100110110111100111101000011001001011101011101111101101110110011000110000101011001001100010100010011111010011010100101100";
	N_in <= "01101010011010101110110010010001111011100111000000110011111111101001001111001101100011000001001000011010011110001011111111110100";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10001011000010111000110100010001011001011001101100111110010010011100110111011100111111011000011000111011110011100110001110110101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01111111100110110111100111101000011001001011101011101111101101110110011000110000101011001001100010100010011111010011010100101100") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=169619234061427452515943317301574317356, exp=56264355201283411649381510693632564085, mod=184822667877625730707730917278973060021";
	REPORT "Expected output is 141453349230748878185067692217169657844, 01101010011010101110110010010001111011100111000000110011111111101001001111001101100011000001001000011010011110001011111111110100";
	N_in <= "01111111100110110111100111101000011001001011101011101111101101110110011000110000101011001001100010100010011111010011010100101100";
	Exp_in <= "00101010010101000001111011100010110011111110101010111101101111010011101100101100011001000011111000000110010111110101101101110101";
	M_in <= "10001011000010111000110100010001011001011001101100111110010010011100110111011100111111011000011000111011110011100110001110110101";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01101010011010101110110010010001111011100111000000110011111111101001001111001101100011000001001000011010011110001011111111110100") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=162011558800030389302711302037615007611, exp=65537, mod=177520508272761769209720826980583177411";
	REPORT "Expected output is 45655028753044940342217127386771013224, 00100010010110001101011010110100111101011101010111001110000101010101100101100010111000001100011101011110100101101011111001101000";
	N_in <= "01111001111000100100101010001110111001100110111111111111101010110100101101000000100010110101110101011111001001011101011101111011";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10000101100011010011010011001101100111110001101111100101101010010111100010100010011111101011000001011010011100010111110011000011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "00100010010110001101011010110100111101011101010111001110000101010101100101100010111000001100011101011110100101101011111001101000") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=45655028753044940342217127386771013224, exp=3602579855696372320547115707745659953, mod=177520508272761769209720826980583177411";
	REPORT "Expected output is 162011558800030389302711302037615007611, 01111001111000100100101010001110111001100110111111111111101010110100101101000000100010110101110101011111001001011101011101111011";
	N_in <= "00100010010110001101011010110100111101011101010111001110000101010101100101100010111000001100011101011110100101101011111001101000";
	Exp_in <= "00000010101101011101010011100110011111110101111000011111100100001101000000101111000111111110101001110000101101110110110000110001";
	M_in <= "10000101100011010011010011001101100111110001101111100101101010010111100010100010011111101011000001011010011100010111110011000011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01111001111000100100101010001110111001100110111111111111101010110100101101000000100010110101110101011111001001011101011101111011") REPORT "test failed" SEVERITY NOTE;


	REPORT "Begin test case for base=156232894051656172687382080664577354971, exp=65537, mod=243815535029074357942427909630916715483";
	REPORT "Expected output is 163821831031182242617884526528449735816, 01111011001111101110111111011110110000010110101111101100110000100101100110011001110101100011010000100011111010111110110010001000";
	N_in <= "01110101100010010101110001100011101000010101010100111010000001110011110011110101011011010101000100100000100010011010110011011011";
	Exp_in <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001";
	M_in <= "10110111011011010010100111111010101110000011110111100111010101000101110000101011101001001011010011000011110110100110001111011011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01111011001111101110111111011110110000010110101111101100110000100101100110011001110101100011010000100011111010111110110010001000") REPORT "test failed" SEVERITY NOTE;

	REPORT "Begin test case for base=163821831031182242617884526528449735816, exp=137356201364243928789970735127789429537, mod=243815535029074357942427909630916715483";
	REPORT "Expected output is 156232894051656172687382080664577354971, 01110101100010010101110001100011101000010101010100111010000001110011110011110101011011010101000100100000100010011010110011011011";
	N_in <= "01111011001111101110111111011110110000010110101111101100110000100101100110011001110101100011010000100011111010111110110010001000";
	Exp_in <= "01100111010101011101011110010101100010001110000001001111000000001010001000001110001001011111110001111101000101011110001100100001";
	M_in <= "10110111011011010010100111111010101110000011110111100111010101000101110000101011101001001011010011000011110110100110001111011011";
	wait for 33409 * clk_period;
	ASSERT(C_out = "01110101100010010101110001100011101000010101010100111010000001110011110011110101011011010101000100100000100010011010110011011011") REPORT "test failed" SEVERITY NOTE;




	wait;

end process;
end;
